
module niosLab2 (
	clk_clk,
	leds_1_name,
	reset_reset_n);	

	input		clk_clk;
	output	[3:0]	leds_1_name;
	input		reset_reset_n;
endmodule
