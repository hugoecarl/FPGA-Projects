// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition"

// DATE "11/12/2020 10:33:45"

// 
// Device: Altera 5CSXFC6D6F31C6 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module niosLab2 (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	clk_clk,
	leds_export,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	clk_clk;
output 	[5:0] leds_export;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \nios2_gen2_0|cpu|W_alu_result[4]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[11]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[10]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[9]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[8]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[7]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[6]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[5]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[12]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[13]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[14]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[15]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[16]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[3]~q ;
wire \nios2_gen2_0|cpu|W_alu_result[2]~q ;
wire \nios2_gen2_0|cpu|F_pc[9]~q ;
wire \nios2_gen2_0|cpu|F_pc[10]~q ;
wire \nios2_gen2_0|cpu|F_pc[11]~q ;
wire \nios2_gen2_0|cpu|F_pc[12]~q ;
wire \nios2_gen2_0|cpu|F_pc[14]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[24] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[25] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[26] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ;
wire \nios2_gen2_0|cpu|F_pc[2]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ;
wire \nios2_gen2_0|cpu|F_pc[8]~q ;
wire \nios2_gen2_0|cpu|F_pc[7]~q ;
wire \nios2_gen2_0|cpu|F_pc[6]~q ;
wire \nios2_gen2_0|cpu|F_pc[5]~q ;
wire \nios2_gen2_0|cpu|F_pc[4]~q ;
wire \nios2_gen2_0|cpu|F_pc[3]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ;
wire \nios2_gen2_0|cpu|F_pc[1]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ;
wire \nios2_gen2_0|cpu|F_pc[0]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[0]~q ;
wire \jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[22]~q ;
wire \nios2_gen2_0|cpu|d_writedata[22]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[23]~q ;
wire \nios2_gen2_0|cpu|d_writedata[23]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[24]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[25]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[26]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[11]~q ;
wire \nios2_gen2_0|cpu|d_writedata[11]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[12]~q ;
wire \nios2_gen2_0|cpu|d_writedata[12]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[13]~q ;
wire \nios2_gen2_0|cpu|d_writedata[13]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[14]~q ;
wire \nios2_gen2_0|cpu|d_writedata[14]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[15]~q ;
wire \nios2_gen2_0|cpu|d_writedata[15]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[16]~q ;
wire \nios2_gen2_0|cpu|d_writedata[16]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[1]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[2]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[3]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[4]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[5]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[8]~q ;
wire \nios2_gen2_0|cpu|d_writedata[8]~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[27] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[28] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[29] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[30] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[31] ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[10]~q ;
wire \nios2_gen2_0|cpu|d_writedata[10]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[17]~q ;
wire \nios2_gen2_0|cpu|d_writedata[17]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[9]~q ;
wire \nios2_gen2_0|cpu|d_writedata[9]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[18]~q ;
wire \nios2_gen2_0|cpu|d_writedata[18]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[19]~q ;
wire \nios2_gen2_0|cpu|d_writedata[19]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[20]~q ;
wire \nios2_gen2_0|cpu|d_writedata[20]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[21]~q ;
wire \nios2_gen2_0|cpu|d_writedata[21]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[16]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[6]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[7]~q ;
wire \jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[27]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[28]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[29]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[30]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[31]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[19]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[18]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[17]~q ;
wire \jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[20]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[21]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[22]~q ;
wire \jtag_uart_0|Add1~1_sumout ;
wire \jtag_uart_0|Add1~5_sumout ;
wire \jtag_uart_0|Add1~9_sumout ;
wire \jtag_uart_0|Add1~13_sumout ;
wire \jtag_uart_0|Add1~17_sumout ;
wire \jtag_uart_0|Add1~21_sumout ;
wire \jtag_uart_0|Add1~25_sumout ;
wire \mm_interconnect_0|nios2_gen2_0_data_master_translator|av_waitrequest~2_combout ;
wire \pio_0|data_out[0]~q ;
wire \pio_0|data_out[1]~q ;
wire \pio_0|data_out[2]~q ;
wire \pio_0|data_out[3]~q ;
wire \pio_0|data_out[4]~q ;
wire \pio_0|data_out[5]~q ;
wire \jtag_uart_0|niosLab2_jtag_uart_0_alt_jtag_atlantic|adapted_tdo~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[0]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|ir_out[0]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|ir_out[1]~q ;
wire \nios2_gen2_0|cpu|d_writedata[0]~q ;
wire \rst_controller|r_sync_rst~q ;
wire \mm_interconnect_0|pio_0_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|router|Equal2~0_combout ;
wire \mm_interconnect_0|router|Equal2~1_combout ;
wire \jtag_uart_0|niosLab2_jtag_uart_0_alt_jtag_atlantic|rst1~q ;
wire \mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[0]~q ;
wire \nios2_gen2_0|cpu|d_write~q ;
wire \mm_interconnect_0|nios2_gen2_0_data_master_translator|write_accepted~q ;
wire \nios2_gen2_0|cpu|d_writedata[1]~q ;
wire \nios2_gen2_0|cpu|d_writedata[2]~q ;
wire \nios2_gen2_0|cpu|d_writedata[3]~q ;
wire \nios2_gen2_0|cpu|d_writedata[4]~q ;
wire \nios2_gen2_0|cpu|d_writedata[5]~q ;
wire \pio_0|always0~3_combout ;
wire \nios2_gen2_0|cpu|d_read~q ;
wire \mm_interconnect_0|nios2_gen2_0_data_master_translator|read_accepted~q ;
wire \jtag_uart_0|always2~0_combout ;
wire \mm_interconnect_0|nios2_gen2_0_data_master_translator|av_waitrequest~0_combout ;
wire \pio_0|always0~4_combout ;
wire \mm_interconnect_0|pio_0_s1_translator|read_latency_shift_reg~1_combout ;
wire \mm_interconnect_0|cmd_mux_001|saved_grant[0]~q ;
wire \nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|waitrequest~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|router|Equal3~0_combout ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \jtag_uart_0|av_waitrequest~q ;
wire \mm_interconnect_0|cmd_demux|WideOr0~3_combout ;
wire \mm_interconnect_0|rsp_demux_002|src0_valid~0_combout ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|rsp_mux|WideOr1~0_combout ;
wire \jtag_uart_0|av_waitrequest~0_combout ;
wire \mm_interconnect_0|cmd_demux|src1_valid~0_combout ;
wire \nios2_gen2_0|cpu|i_read~q ;
wire \nios2_gen2_0|cpu|F_pc[13]~q ;
wire \mm_interconnect_0|cmd_mux_001|src_valid~0_combout ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem~0_combout ;
wire \mm_interconnect_0|cmd_demux|src2_valid~0_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_valid~0_combout ;
wire \nios2_gen2_0|cpu|hbreak_enabled~q ;
wire \mm_interconnect_0|nios2_gen2_0_data_master_translator|av_waitrequest~1_combout ;
wire \mm_interconnect_0|rsp_demux_001|src0_valid~0_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[0]~combout ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[22]~q ;
wire \mm_interconnect_0|rsp_demux_001|src1_valid~0_combout ;
wire \mm_interconnect_0|rsp_demux_002|src1_valid~0_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[22]~combout ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[23]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_data[23]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[24]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[25]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[26]~combout ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[11]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[12]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_data[12]~combout ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[13]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[14]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_data[14]~combout ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[15]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[16]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_data[0]~combout ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[1]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_data[2]~combout ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[3]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[4]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[5]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[8]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_data[8]~combout ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[10]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_data[10]~combout ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[17]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_data[17]~combout ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[9]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_data[9]~combout ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[18]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[19]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[20]~q ;
wire \mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[21]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_data[6]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[46]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[7]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[1]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[2]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[3]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[4]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[5]~combout ;
wire \jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \rst_controller|r_early_rst~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[46]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[47]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[48]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[49]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[50]~combout ;
wire \nios2_gen2_0|cpu|d_byteenable[0]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[32]~combout ;
wire \jtag_uart_0|ien_AF~q ;
wire \jtag_uart_0|read_0~q ;
wire \pio_0|readdata[0]~0_combout ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[8]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~1_combout ;
wire \nios2_gen2_0|cpu|d_byteenable[2]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[34]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~2_combout ;
wire \nios2_gen2_0|cpu|d_writedata[24]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~3_combout ;
wire \nios2_gen2_0|cpu|d_byteenable[3]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[35]~combout ;
wire \nios2_gen2_0|cpu|d_writedata[25]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~4_combout ;
wire \nios2_gen2_0|cpu|d_writedata[26]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~5_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~6_combout ;
wire \nios2_gen2_0|cpu|d_byteenable[1]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[33]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~17_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[27]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[28]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[29]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[30]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[31]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~19_combout ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[10]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[9]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~0_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~1_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~20_combout ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[12]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~21_combout ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[13]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~22_combout ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[14]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~23_combout ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[15]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~24_combout ;
wire \nios2_gen2_0|cpu|d_writedata[6]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~25_combout ;
wire \nios2_gen2_0|cpu|d_writedata[7]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~26_combout ;
wire \jtag_uart_0|ien_AE~q ;
wire \pio_0|readdata[1]~1_combout ;
wire \pio_0|readdata[2]~2_combout ;
wire \pio_0|readdata[3]~3_combout ;
wire \pio_0|readdata[4]~4_combout ;
wire \pio_0|readdata[5]~5_combout ;
wire \jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~1_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[32]~combout ;
wire \jtag_uart_0|av_readdata[8]~0_combout ;
wire \nios2_gen2_0|cpu|d_writedata[27]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~27_combout ;
wire \nios2_gen2_0|cpu|d_writedata[28]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~28_combout ;
wire \nios2_gen2_0|cpu|d_writedata[29]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~29_combout ;
wire \nios2_gen2_0|cpu|d_writedata[30]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~30_combout ;
wire \nios2_gen2_0|cpu|d_writedata[31]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~31_combout ;
wire \jtag_uart_0|ac~q ;
wire \jtag_uart_0|av_readdata[9]~combout ;
wire \jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \jtag_uart_0|woverflow~q ;
wire \jtag_uart_0|rvalid~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~2_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~2_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~3_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~4_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~5_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~6_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~7_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~8_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~3_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~4_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~5_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[34]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[35]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[33]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~19_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~20_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~22_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~23_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~24_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~25_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~26_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~27_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~28_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~29_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~30_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~31_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~32_combout ;
wire \rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ;
wire \~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \clk_clk~input_o ;
wire \reset_reset_n~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \altera_internal_jtag~TDIUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \altera_internal_jtag~TDO ;


niosLab2_altera_reset_controller rst_controller(
	.r_sync_rst1(\rst_controller|r_sync_rst~q ),
	.r_early_rst1(\rst_controller|r_early_rst~q ),
	.altera_reset_synchronizer_int_chain_1(\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

niosLab2_niosLab2_nios2_gen2_0 nios2_gen2_0(
	.W_alu_result_4(\nios2_gen2_0|cpu|W_alu_result[4]~q ),
	.W_alu_result_11(\nios2_gen2_0|cpu|W_alu_result[11]~q ),
	.W_alu_result_10(\nios2_gen2_0|cpu|W_alu_result[10]~q ),
	.W_alu_result_9(\nios2_gen2_0|cpu|W_alu_result[9]~q ),
	.W_alu_result_8(\nios2_gen2_0|cpu|W_alu_result[8]~q ),
	.W_alu_result_7(\nios2_gen2_0|cpu|W_alu_result[7]~q ),
	.W_alu_result_6(\nios2_gen2_0|cpu|W_alu_result[6]~q ),
	.W_alu_result_5(\nios2_gen2_0|cpu|W_alu_result[5]~q ),
	.W_alu_result_12(\nios2_gen2_0|cpu|W_alu_result[12]~q ),
	.W_alu_result_13(\nios2_gen2_0|cpu|W_alu_result[13]~q ),
	.W_alu_result_14(\nios2_gen2_0|cpu|W_alu_result[14]~q ),
	.W_alu_result_15(\nios2_gen2_0|cpu|W_alu_result[15]~q ),
	.W_alu_result_16(\nios2_gen2_0|cpu|W_alu_result[16]~q ),
	.W_alu_result_3(\nios2_gen2_0|cpu|W_alu_result[3]~q ),
	.W_alu_result_2(\nios2_gen2_0|cpu|W_alu_result[2]~q ),
	.F_pc_9(\nios2_gen2_0|cpu|F_pc[9]~q ),
	.F_pc_10(\nios2_gen2_0|cpu|F_pc[10]~q ),
	.F_pc_11(\nios2_gen2_0|cpu|F_pc[11]~q ),
	.F_pc_12(\nios2_gen2_0|cpu|F_pc[12]~q ),
	.F_pc_14(\nios2_gen2_0|cpu|F_pc[14]~q ),
	.q_a_22(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_23(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_11(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_12(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_13(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_14(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_15(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_16(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_1(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_3(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_4(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_5(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ),
	.F_pc_2(\nios2_gen2_0|cpu|F_pc[2]~q ),
	.q_a_8(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_10(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_17(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ),
	.F_pc_8(\nios2_gen2_0|cpu|F_pc[8]~q ),
	.F_pc_7(\nios2_gen2_0|cpu|F_pc[7]~q ),
	.F_pc_6(\nios2_gen2_0|cpu|F_pc[6]~q ),
	.F_pc_5(\nios2_gen2_0|cpu|F_pc[5]~q ),
	.F_pc_4(\nios2_gen2_0|cpu|F_pc[4]~q ),
	.F_pc_3(\nios2_gen2_0|cpu|F_pc[3]~q ),
	.q_a_9(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_18(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_19(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_20(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_21(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ),
	.F_pc_1(\nios2_gen2_0|cpu|F_pc[1]~q ),
	.F_pc_0(\nios2_gen2_0|cpu|F_pc[0]~q ),
	.readdata_0(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[0]~q ),
	.readdata_22(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[22]~q ),
	.d_writedata_22(\nios2_gen2_0|cpu|d_writedata[22]~q ),
	.readdata_23(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[23]~q ),
	.d_writedata_23(\nios2_gen2_0|cpu|d_writedata[23]~q ),
	.readdata_24(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[24]~q ),
	.readdata_25(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[25]~q ),
	.readdata_26(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[26]~q ),
	.readdata_11(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[11]~q ),
	.d_writedata_11(\nios2_gen2_0|cpu|d_writedata[11]~q ),
	.readdata_12(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[12]~q ),
	.d_writedata_12(\nios2_gen2_0|cpu|d_writedata[12]~q ),
	.readdata_13(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[13]~q ),
	.d_writedata_13(\nios2_gen2_0|cpu|d_writedata[13]~q ),
	.readdata_14(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[14]~q ),
	.d_writedata_14(\nios2_gen2_0|cpu|d_writedata[14]~q ),
	.readdata_15(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[15]~q ),
	.d_writedata_15(\nios2_gen2_0|cpu|d_writedata[15]~q ),
	.readdata_16(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[16]~q ),
	.d_writedata_16(\nios2_gen2_0|cpu|d_writedata[16]~q ),
	.readdata_1(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[1]~q ),
	.readdata_2(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[2]~q ),
	.readdata_3(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[3]~q ),
	.readdata_4(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[4]~q ),
	.readdata_5(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[5]~q ),
	.readdata_8(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[8]~q ),
	.d_writedata_8(\nios2_gen2_0|cpu|d_writedata[8]~q ),
	.readdata_10(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[10]~q ),
	.d_writedata_10(\nios2_gen2_0|cpu|d_writedata[10]~q ),
	.readdata_17(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[17]~q ),
	.d_writedata_17(\nios2_gen2_0|cpu|d_writedata[17]~q ),
	.readdata_9(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[9]~q ),
	.d_writedata_9(\nios2_gen2_0|cpu|d_writedata[9]~q ),
	.readdata_18(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[18]~q ),
	.d_writedata_18(\nios2_gen2_0|cpu|d_writedata[18]~q ),
	.readdata_19(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[19]~q ),
	.d_writedata_19(\nios2_gen2_0|cpu|d_writedata[19]~q ),
	.readdata_20(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[20]~q ),
	.d_writedata_20(\nios2_gen2_0|cpu|d_writedata[20]~q ),
	.readdata_21(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[21]~q ),
	.d_writedata_21(\nios2_gen2_0|cpu|d_writedata[21]~q ),
	.av_readdata_pre_16(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.readdata_6(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[6]~q ),
	.readdata_7(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[7]~q ),
	.readdata_27(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[27]~q ),
	.readdata_28(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[28]~q ),
	.readdata_29(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[29]~q ),
	.readdata_30(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[30]~q ),
	.readdata_31(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[31]~q ),
	.av_readdata_pre_19(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_18(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_17(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_20(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_21(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_22(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.av_waitrequest(\mm_interconnect_0|nios2_gen2_0_data_master_translator|av_waitrequest~2_combout ),
	.sr_0(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[0]~q ),
	.ir_out_0(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|ir_out[0]~q ),
	.ir_out_1(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|ir_out[1]~q ),
	.d_writedata_0(\nios2_gen2_0|cpu|d_writedata[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.d_write(\nios2_gen2_0|cpu|d_write~q ),
	.d_writedata_1(\nios2_gen2_0|cpu|d_writedata[1]~q ),
	.d_writedata_2(\nios2_gen2_0|cpu|d_writedata[2]~q ),
	.d_writedata_3(\nios2_gen2_0|cpu|d_writedata[3]~q ),
	.d_writedata_4(\nios2_gen2_0|cpu|d_writedata[4]~q ),
	.d_writedata_5(\nios2_gen2_0|cpu|d_writedata[5]~q ),
	.d_read(\nios2_gen2_0|cpu|d_read~q ),
	.always2(\jtag_uart_0|always2~0_combout ),
	.av_waitrequest1(\mm_interconnect_0|nios2_gen2_0_data_master_translator|av_waitrequest~0_combout ),
	.read_latency_shift_reg(\mm_interconnect_0|pio_0_s1_translator|read_latency_shift_reg~1_combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_001|saved_grant[0]~q ),
	.debug_mem_slave_waitrequest(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\mm_interconnect_0|cmd_demux|WideOr0~3_combout ),
	.src0_valid(\mm_interconnect_0|rsp_demux_002|src0_valid~0_combout ),
	.read_latency_shift_reg_0(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~0_combout ),
	.src1_valid(\mm_interconnect_0|cmd_demux|src1_valid~0_combout ),
	.i_read(\nios2_gen2_0|cpu|i_read~q ),
	.F_pc_13(\nios2_gen2_0|cpu|F_pc[13]~q ),
	.src_valid(\mm_interconnect_0|cmd_mux_001|src_valid~0_combout ),
	.mem(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem~0_combout ),
	.hbreak_enabled(\nios2_gen2_0|cpu|hbreak_enabled~q ),
	.av_waitrequest2(\mm_interconnect_0|nios2_gen2_0_data_master_translator|av_waitrequest~1_combout ),
	.src0_valid1(\mm_interconnect_0|rsp_demux_001|src0_valid~0_combout ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~combout ),
	.av_readdata_pre_221(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[22]~q ),
	.src1_valid1(\mm_interconnect_0|rsp_demux_001|src1_valid~0_combout ),
	.src1_valid2(\mm_interconnect_0|rsp_demux_002|src1_valid~0_combout ),
	.src_data_22(\mm_interconnect_0|rsp_mux_001|src_data[22]~combout ),
	.av_readdata_pre_23(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[23]~q ),
	.src_data_23(\mm_interconnect_0|rsp_mux_001|src_data[23]~combout ),
	.src_data_24(\mm_interconnect_0|rsp_mux_001|src_data[24]~combout ),
	.src_data_25(\mm_interconnect_0|rsp_mux_001|src_data[25]~combout ),
	.src_data_26(\mm_interconnect_0|rsp_mux_001|src_data[26]~combout ),
	.av_readdata_pre_11(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_12(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[12]~q ),
	.src_data_12(\mm_interconnect_0|rsp_mux_001|src_data[12]~combout ),
	.av_readdata_pre_13(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[14]~q ),
	.src_data_14(\mm_interconnect_0|rsp_mux_001|src_data[14]~combout ),
	.av_readdata_pre_15(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_161(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[16]~q ),
	.src_data_01(\mm_interconnect_0|rsp_mux_001|src_data[0]~combout ),
	.av_readdata_pre_1(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[1]~q ),
	.src_data_2(\mm_interconnect_0|rsp_mux_001|src_data[2]~combout ),
	.av_readdata_pre_3(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_8(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[8]~q ),
	.src_data_8(\mm_interconnect_0|rsp_mux_001|src_data[8]~combout ),
	.av_readdata_pre_10(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[10]~q ),
	.src_data_10(\mm_interconnect_0|rsp_mux_001|src_data[10]~combout ),
	.av_readdata_pre_171(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[17]~q ),
	.src_data_17(\mm_interconnect_0|rsp_mux_001|src_data[17]~combout ),
	.av_readdata_pre_9(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[9]~q ),
	.src_data_9(\mm_interconnect_0|rsp_mux_001|src_data[9]~combout ),
	.av_readdata_pre_181(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_191(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_201(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_211(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[21]~q ),
	.src_data_6(\mm_interconnect_0|rsp_mux_001|src_data[6]~combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_001|src_data[46]~combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux_001|src_data[7]~combout ),
	.src_data_1(\mm_interconnect_0|rsp_mux|src_data[1]~combout ),
	.src_data_21(\mm_interconnect_0|rsp_mux|src_data[2]~combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux|src_data[3]~combout ),
	.src_data_4(\mm_interconnect_0|rsp_mux|src_data[4]~combout ),
	.src_data_5(\mm_interconnect_0|rsp_mux|src_data[5]~combout ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.d_byteenable_0(\nios2_gen2_0|cpu|d_byteenable[0]~q ),
	.av_readdata_pre_81(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.d_byteenable_2(\nios2_gen2_0|cpu|d_byteenable[2]~q ),
	.d_writedata_24(\nios2_gen2_0|cpu|d_writedata[24]~q ),
	.d_byteenable_3(\nios2_gen2_0|cpu|d_byteenable[3]~q ),
	.d_writedata_25(\nios2_gen2_0|cpu|d_writedata[25]~q ),
	.d_writedata_26(\nios2_gen2_0|cpu|d_writedata[26]~q ),
	.d_byteenable_1(\nios2_gen2_0|cpu|d_byteenable[1]~q ),
	.src_data_27(\mm_interconnect_0|rsp_mux_001|src_data[27]~combout ),
	.src_data_28(\mm_interconnect_0|rsp_mux_001|src_data[28]~combout ),
	.src_data_29(\mm_interconnect_0|rsp_mux_001|src_data[29]~combout ),
	.src_data_30(\mm_interconnect_0|rsp_mux_001|src_data[30]~combout ),
	.src_data_31(\mm_interconnect_0|rsp_mux_001|src_data[31]~combout ),
	.av_readdata_pre_101(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_91(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.src_payload(\mm_interconnect_0|rsp_mux|src_payload~0_combout ),
	.src_payload1(\mm_interconnect_0|rsp_mux|src_payload~1_combout ),
	.av_readdata_pre_121(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_131(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_141(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_151(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.d_writedata_6(\nios2_gen2_0|cpu|d_writedata[6]~q ),
	.d_writedata_7(\nios2_gen2_0|cpu|d_writedata[7]~q ),
	.src_payload2(\mm_interconnect_0|cmd_mux_001|src_payload~0_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_001|src_data[38]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_001|src_data[41]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_001|src_data[45]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_001|src_data[44]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_001|src_data[43]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_001|src_data[42]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_001|src_data[40]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_001|src_data[39]~combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_001|src_payload~1_combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_001|src_data[32]~combout ),
	.d_writedata_27(\nios2_gen2_0|cpu|d_writedata[27]~q ),
	.d_writedata_28(\nios2_gen2_0|cpu|d_writedata[28]~q ),
	.d_writedata_29(\nios2_gen2_0|cpu|d_writedata[29]~q ),
	.d_writedata_30(\nios2_gen2_0|cpu|d_writedata[30]~q ),
	.d_writedata_31(\nios2_gen2_0|cpu|d_writedata[31]~q ),
	.src_payload4(\mm_interconnect_0|rsp_mux|src_payload~2_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_001|src_payload~2_combout ),
	.src_payload6(\mm_interconnect_0|rsp_mux|src_payload~3_combout ),
	.src_payload7(\mm_interconnect_0|rsp_mux|src_payload~4_combout ),
	.src_payload8(\mm_interconnect_0|rsp_mux|src_payload~5_combout ),
	.src_payload9(\mm_interconnect_0|rsp_mux|src_payload~6_combout ),
	.src_payload10(\mm_interconnect_0|rsp_mux|src_payload~7_combout ),
	.src_payload11(\mm_interconnect_0|rsp_mux|src_payload~8_combout ),
	.src_payload12(\mm_interconnect_0|rsp_mux|src_payload~9_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_001|src_payload~3_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_001|src_payload~4_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_001|src_payload~5_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_001|src_data[34]~combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_001|src_payload~6_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_001|src_payload~7_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_001|src_data[35]~combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_001|src_payload~8_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_001|src_payload~9_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_001|src_payload~10_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_001|src_data[33]~combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_001|src_payload~11_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_001|src_payload~12_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_001|src_payload~13_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_001|src_payload~14_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_001|src_payload~15_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_001|src_payload~16_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_001|src_payload~17_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_001|src_payload~18_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_001|src_payload~19_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_001|src_payload~20_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_001|src_payload~21_combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_001|src_payload~22_combout ),
	.src_payload33(\mm_interconnect_0|cmd_mux_001|src_payload~23_combout ),
	.src_payload34(\mm_interconnect_0|cmd_mux_001|src_payload~24_combout ),
	.src_payload35(\mm_interconnect_0|cmd_mux_001|src_payload~25_combout ),
	.src_payload36(\mm_interconnect_0|cmd_mux_001|src_payload~26_combout ),
	.src_payload37(\mm_interconnect_0|cmd_mux_001|src_payload~27_combout ),
	.src_payload38(\mm_interconnect_0|cmd_mux_001|src_payload~28_combout ),
	.src_payload39(\mm_interconnect_0|cmd_mux_001|src_payload~29_combout ),
	.src_payload40(\mm_interconnect_0|cmd_mux_001|src_payload~30_combout ),
	.src_payload41(\mm_interconnect_0|cmd_mux_001|src_payload~31_combout ),
	.src_payload42(\mm_interconnect_0|cmd_mux_001|src_payload~32_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.splitter_nodes_receive_1_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.irf_reg_0_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.irf_reg_1_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.clk_clk(\clk_clk~input_o ));

niosLab2_niosLab2_mm_interconnect_0 mm_interconnect_0(
	.W_alu_result_4(\nios2_gen2_0|cpu|W_alu_result[4]~q ),
	.W_alu_result_11(\nios2_gen2_0|cpu|W_alu_result[11]~q ),
	.W_alu_result_10(\nios2_gen2_0|cpu|W_alu_result[10]~q ),
	.W_alu_result_9(\nios2_gen2_0|cpu|W_alu_result[9]~q ),
	.W_alu_result_8(\nios2_gen2_0|cpu|W_alu_result[8]~q ),
	.W_alu_result_7(\nios2_gen2_0|cpu|W_alu_result[7]~q ),
	.W_alu_result_6(\nios2_gen2_0|cpu|W_alu_result[6]~q ),
	.W_alu_result_5(\nios2_gen2_0|cpu|W_alu_result[5]~q ),
	.W_alu_result_12(\nios2_gen2_0|cpu|W_alu_result[12]~q ),
	.W_alu_result_13(\nios2_gen2_0|cpu|W_alu_result[13]~q ),
	.W_alu_result_14(\nios2_gen2_0|cpu|W_alu_result[14]~q ),
	.W_alu_result_15(\nios2_gen2_0|cpu|W_alu_result[15]~q ),
	.W_alu_result_16(\nios2_gen2_0|cpu|W_alu_result[16]~q ),
	.W_alu_result_3(\nios2_gen2_0|cpu|W_alu_result[3]~q ),
	.W_alu_result_2(\nios2_gen2_0|cpu|W_alu_result[2]~q ),
	.F_pc_9(\nios2_gen2_0|cpu|F_pc[9]~q ),
	.F_pc_10(\nios2_gen2_0|cpu|F_pc[10]~q ),
	.F_pc_11(\nios2_gen2_0|cpu|F_pc[11]~q ),
	.F_pc_12(\nios2_gen2_0|cpu|F_pc[12]~q ),
	.F_pc_14(\nios2_gen2_0|cpu|F_pc[14]~q ),
	.q_a_0(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_22(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_23(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_24(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_25(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_26(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_12(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_14(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_1(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_2(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_3(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_4(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_5(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ),
	.F_pc_2(\nios2_gen2_0|cpu|F_pc[2]~q ),
	.q_a_8(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_10(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_17(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ),
	.F_pc_8(\nios2_gen2_0|cpu|F_pc[8]~q ),
	.F_pc_7(\nios2_gen2_0|cpu|F_pc[7]~q ),
	.F_pc_6(\nios2_gen2_0|cpu|F_pc[6]~q ),
	.F_pc_5(\nios2_gen2_0|cpu|F_pc[5]~q ),
	.F_pc_4(\nios2_gen2_0|cpu|F_pc[4]~q ),
	.F_pc_3(\nios2_gen2_0|cpu|F_pc[3]~q ),
	.q_a_9(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_6(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ),
	.F_pc_1(\nios2_gen2_0|cpu|F_pc[1]~q ),
	.q_a_7(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ),
	.F_pc_0(\nios2_gen2_0|cpu|F_pc[0]~q ),
	.readdata_0(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[0]~q ),
	.q_b_0(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.readdata_22(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[22]~q ),
	.d_writedata_22(\nios2_gen2_0|cpu|d_writedata[22]~q ),
	.readdata_23(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[23]~q ),
	.d_writedata_23(\nios2_gen2_0|cpu|d_writedata[23]~q ),
	.readdata_24(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[24]~q ),
	.readdata_25(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[25]~q ),
	.readdata_26(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[26]~q ),
	.readdata_11(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[11]~q ),
	.d_writedata_11(\nios2_gen2_0|cpu|d_writedata[11]~q ),
	.readdata_12(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[12]~q ),
	.d_writedata_12(\nios2_gen2_0|cpu|d_writedata[12]~q ),
	.readdata_13(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[13]~q ),
	.d_writedata_13(\nios2_gen2_0|cpu|d_writedata[13]~q ),
	.readdata_14(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[14]~q ),
	.d_writedata_14(\nios2_gen2_0|cpu|d_writedata[14]~q ),
	.readdata_15(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[15]~q ),
	.d_writedata_15(\nios2_gen2_0|cpu|d_writedata[15]~q ),
	.readdata_16(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[16]~q ),
	.d_writedata_16(\nios2_gen2_0|cpu|d_writedata[16]~q ),
	.readdata_1(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[1]~q ),
	.readdata_2(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[2]~q ),
	.readdata_3(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[3]~q ),
	.readdata_4(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[4]~q ),
	.readdata_5(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[5]~q ),
	.readdata_8(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[8]~q ),
	.d_writedata_8(\nios2_gen2_0|cpu|d_writedata[8]~q ),
	.q_a_27(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_28(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_29(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_30(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_31(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[31] ),
	.readdata_10(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[10]~q ),
	.d_writedata_10(\nios2_gen2_0|cpu|d_writedata[10]~q ),
	.readdata_17(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[17]~q ),
	.d_writedata_17(\nios2_gen2_0|cpu|d_writedata[17]~q ),
	.readdata_9(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[9]~q ),
	.d_writedata_9(\nios2_gen2_0|cpu|d_writedata[9]~q ),
	.readdata_18(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[18]~q ),
	.d_writedata_18(\nios2_gen2_0|cpu|d_writedata[18]~q ),
	.readdata_19(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[19]~q ),
	.d_writedata_19(\nios2_gen2_0|cpu|d_writedata[19]~q ),
	.readdata_20(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[20]~q ),
	.d_writedata_20(\nios2_gen2_0|cpu|d_writedata[20]~q ),
	.readdata_21(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[21]~q ),
	.d_writedata_21(\nios2_gen2_0|cpu|d_writedata[21]~q ),
	.av_readdata_pre_16(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.readdata_6(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[6]~q ),
	.readdata_7(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[7]~q ),
	.q_b_1(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.readdata_27(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[27]~q ),
	.readdata_28(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[28]~q ),
	.readdata_29(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[29]~q ),
	.readdata_30(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[30]~q ),
	.readdata_31(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|readdata[31]~q ),
	.av_readdata_pre_19(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_18(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_17(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.q_b_7(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_6(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.av_readdata_pre_20(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_21(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_22(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.Add1(\jtag_uart_0|Add1~1_sumout ),
	.Add11(\jtag_uart_0|Add1~5_sumout ),
	.Add12(\jtag_uart_0|Add1~9_sumout ),
	.Add13(\jtag_uart_0|Add1~13_sumout ),
	.Add14(\jtag_uart_0|Add1~17_sumout ),
	.Add15(\jtag_uart_0|Add1~21_sumout ),
	.Add16(\jtag_uart_0|Add1~25_sumout ),
	.nios2_gen2_0_data_master_waitrequest(\mm_interconnect_0|nios2_gen2_0_data_master_translator|av_waitrequest~2_combout ),
	.d_writedata_0(\nios2_gen2_0|cpu|d_writedata[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.mem_used_1(\mm_interconnect_0|pio_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.Equal2(\mm_interconnect_0|router|Equal2~0_combout ),
	.Equal21(\mm_interconnect_0|router|Equal2~1_combout ),
	.rst1(\jtag_uart_0|niosLab2_jtag_uart_0_alt_jtag_atlantic|rst1~q ),
	.wait_latency_counter_1(\mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[0]~q ),
	.d_write(\nios2_gen2_0|cpu|d_write~q ),
	.write_accepted(\mm_interconnect_0|nios2_gen2_0_data_master_translator|write_accepted~q ),
	.d_writedata_1(\nios2_gen2_0|cpu|d_writedata[1]~q ),
	.d_writedata_2(\nios2_gen2_0|cpu|d_writedata[2]~q ),
	.d_writedata_3(\nios2_gen2_0|cpu|d_writedata[3]~q ),
	.d_writedata_4(\nios2_gen2_0|cpu|d_writedata[4]~q ),
	.d_writedata_5(\nios2_gen2_0|cpu|d_writedata[5]~q ),
	.always0(\pio_0|always0~3_combout ),
	.d_read(\nios2_gen2_0|cpu|d_read~q ),
	.read_accepted(\mm_interconnect_0|nios2_gen2_0_data_master_translator|read_accepted~q ),
	.always2(\jtag_uart_0|always2~0_combout ),
	.av_waitrequest(\mm_interconnect_0|nios2_gen2_0_data_master_translator|av_waitrequest~0_combout ),
	.always01(\pio_0|always0~4_combout ),
	.read_latency_shift_reg(\mm_interconnect_0|pio_0_s1_translator|read_latency_shift_reg~1_combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_001|saved_grant[0]~q ),
	.waitrequest(\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|waitrequest~q ),
	.mem_used_11(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ),
	.saved_grant_01(\mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ),
	.mem_used_12(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.Equal3(\mm_interconnect_0|router|Equal3~0_combout ),
	.mem_used_13(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest1(\jtag_uart_0|av_waitrequest~q ),
	.WideOr0(\mm_interconnect_0|cmd_demux|WideOr0~3_combout ),
	.src0_valid(\mm_interconnect_0|rsp_demux_002|src0_valid~0_combout ),
	.read_latency_shift_reg_0(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~0_combout ),
	.av_waitrequest2(\jtag_uart_0|av_waitrequest~0_combout ),
	.src1_valid(\mm_interconnect_0|cmd_demux|src1_valid~0_combout ),
	.i_read(\nios2_gen2_0|cpu|i_read~q ),
	.F_pc_13(\nios2_gen2_0|cpu|F_pc[13]~q ),
	.src_valid(\mm_interconnect_0|cmd_mux_001|src_valid~0_combout ),
	.mem(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem~0_combout ),
	.src2_valid(\mm_interconnect_0|cmd_demux|src2_valid~0_combout ),
	.src_valid1(\mm_interconnect_0|cmd_mux_002|src_valid~0_combout ),
	.hbreak_enabled(\nios2_gen2_0|cpu|hbreak_enabled~q ),
	.av_waitrequest3(\mm_interconnect_0|nios2_gen2_0_data_master_translator|av_waitrequest~1_combout ),
	.src0_valid1(\mm_interconnect_0|rsp_demux_001|src0_valid~0_combout ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~combout ),
	.av_readdata_pre_221(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[22]~q ),
	.src1_valid1(\mm_interconnect_0|rsp_demux_001|src1_valid~0_combout ),
	.src1_valid2(\mm_interconnect_0|rsp_demux_002|src1_valid~0_combout ),
	.src_data_22(\mm_interconnect_0|rsp_mux_001|src_data[22]~combout ),
	.av_readdata_pre_23(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[23]~q ),
	.src_data_23(\mm_interconnect_0|rsp_mux_001|src_data[23]~combout ),
	.src_data_24(\mm_interconnect_0|rsp_mux_001|src_data[24]~combout ),
	.src_data_25(\mm_interconnect_0|rsp_mux_001|src_data[25]~combout ),
	.src_data_26(\mm_interconnect_0|rsp_mux_001|src_data[26]~combout ),
	.av_readdata_pre_11(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_12(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[12]~q ),
	.src_data_12(\mm_interconnect_0|rsp_mux_001|src_data[12]~combout ),
	.av_readdata_pre_13(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[14]~q ),
	.src_data_14(\mm_interconnect_0|rsp_mux_001|src_data[14]~combout ),
	.av_readdata_pre_15(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_161(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[16]~q ),
	.src_data_01(\mm_interconnect_0|rsp_mux_001|src_data[0]~combout ),
	.av_readdata_pre_1(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[1]~q ),
	.src_data_2(\mm_interconnect_0|rsp_mux_001|src_data[2]~combout ),
	.av_readdata_pre_3(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_8(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[8]~q ),
	.src_data_8(\mm_interconnect_0|rsp_mux_001|src_data[8]~combout ),
	.av_readdata_pre_10(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[10]~q ),
	.src_data_10(\mm_interconnect_0|rsp_mux_001|src_data[10]~combout ),
	.av_readdata_pre_171(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[17]~q ),
	.src_data_17(\mm_interconnect_0|rsp_mux_001|src_data[17]~combout ),
	.av_readdata_pre_9(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[9]~q ),
	.src_data_9(\mm_interconnect_0|rsp_mux_001|src_data[9]~combout ),
	.av_readdata_pre_181(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_191(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_201(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_211(\mm_interconnect_0|nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[21]~q ),
	.src_data_6(\mm_interconnect_0|rsp_mux_001|src_data[6]~combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_001|src_data[46]~combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux_001|src_data[7]~combout ),
	.src_data_1(\mm_interconnect_0|rsp_mux|src_data[1]~combout ),
	.src_data_21(\mm_interconnect_0|rsp_mux|src_data[2]~combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux|src_data[3]~combout ),
	.src_data_4(\mm_interconnect_0|rsp_mux|src_data[4]~combout ),
	.src_data_5(\mm_interconnect_0|rsp_mux|src_data[5]~combout ),
	.b_full(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_002|src_payload~0_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_002|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_002|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_002|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_002|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_002|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_002|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_002|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_002|src_data[45]~combout ),
	.src_data_461(\mm_interconnect_0|cmd_mux_002|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_0|cmd_mux_002|src_data[47]~combout ),
	.src_data_48(\mm_interconnect_0|cmd_mux_002|src_data[48]~combout ),
	.src_data_49(\mm_interconnect_0|cmd_mux_002|src_data[49]~combout ),
	.src_data_50(\mm_interconnect_0|cmd_mux_002|src_data[50]~combout ),
	.d_byteenable_0(\nios2_gen2_0|cpu|d_byteenable[0]~q ),
	.src_data_32(\mm_interconnect_0|cmd_mux_002|src_data[32]~combout ),
	.ien_AF(\jtag_uart_0|ien_AF~q ),
	.read_0(\jtag_uart_0|read_0~q ),
	.readdata_01(\pio_0|readdata[0]~0_combout ),
	.av_readdata_pre_81(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.src_payload1(\mm_interconnect_0|cmd_mux_002|src_payload~1_combout ),
	.d_byteenable_2(\nios2_gen2_0|cpu|d_byteenable[2]~q ),
	.src_data_34(\mm_interconnect_0|cmd_mux_002|src_data[34]~combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_002|src_payload~2_combout ),
	.d_writedata_24(\nios2_gen2_0|cpu|d_writedata[24]~q ),
	.src_payload3(\mm_interconnect_0|cmd_mux_002|src_payload~3_combout ),
	.d_byteenable_3(\nios2_gen2_0|cpu|d_byteenable[3]~q ),
	.src_data_35(\mm_interconnect_0|cmd_mux_002|src_data[35]~combout ),
	.d_writedata_25(\nios2_gen2_0|cpu|d_writedata[25]~q ),
	.src_payload4(\mm_interconnect_0|cmd_mux_002|src_payload~4_combout ),
	.d_writedata_26(\nios2_gen2_0|cpu|d_writedata[26]~q ),
	.src_payload5(\mm_interconnect_0|cmd_mux_002|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_002|src_payload~6_combout ),
	.d_byteenable_1(\nios2_gen2_0|cpu|d_byteenable[1]~q ),
	.src_data_33(\mm_interconnect_0|cmd_mux_002|src_data[33]~combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_002|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_002|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_002|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_002|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_002|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_002|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_002|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_002|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_002|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_002|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_002|src_payload~17_combout ),
	.src_data_27(\mm_interconnect_0|rsp_mux_001|src_data[27]~combout ),
	.src_data_28(\mm_interconnect_0|rsp_mux_001|src_data[28]~combout ),
	.src_data_29(\mm_interconnect_0|rsp_mux_001|src_data[29]~combout ),
	.src_data_30(\mm_interconnect_0|rsp_mux_001|src_data[30]~combout ),
	.src_data_31(\mm_interconnect_0|rsp_mux_001|src_data[31]~combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_002|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_002|src_payload~19_combout ),
	.av_readdata_pre_101(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_91(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.src_payload20(\mm_interconnect_0|rsp_mux|src_payload~0_combout ),
	.src_payload21(\mm_interconnect_0|rsp_mux|src_payload~1_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_002|src_payload~20_combout ),
	.av_readdata_pre_121(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.src_payload23(\mm_interconnect_0|cmd_mux_002|src_payload~21_combout ),
	.av_readdata_pre_131(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.src_payload24(\mm_interconnect_0|cmd_mux_002|src_payload~22_combout ),
	.av_readdata_pre_141(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.src_payload25(\mm_interconnect_0|cmd_mux_002|src_payload~23_combout ),
	.av_readdata_pre_151(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.src_payload26(\mm_interconnect_0|cmd_mux_002|src_payload~24_combout ),
	.d_writedata_6(\nios2_gen2_0|cpu|d_writedata[6]~q ),
	.src_payload27(\mm_interconnect_0|cmd_mux_002|src_payload~25_combout ),
	.d_writedata_7(\nios2_gen2_0|cpu|d_writedata[7]~q ),
	.src_payload28(\mm_interconnect_0|cmd_mux_002|src_payload~26_combout ),
	.ien_AE(\jtag_uart_0|ien_AE~q ),
	.readdata_110(\pio_0|readdata[1]~1_combout ),
	.readdata_210(\pio_0|readdata[2]~2_combout ),
	.readdata_32(\pio_0|readdata[3]~3_combout ),
	.readdata_41(\pio_0|readdata[4]~4_combout ),
	.readdata_51(\pio_0|readdata[5]~5_combout ),
	.b_non_empty(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.counter_reg_bit_1(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_5(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.src_payload29(\mm_interconnect_0|cmd_mux_001|src_payload~0_combout ),
	.src_data_381(\mm_interconnect_0|cmd_mux_001|src_data[38]~combout ),
	.src_data_411(\mm_interconnect_0|cmd_mux_001|src_data[41]~combout ),
	.src_data_451(\mm_interconnect_0|cmd_mux_001|src_data[45]~combout ),
	.src_data_441(\mm_interconnect_0|cmd_mux_001|src_data[44]~combout ),
	.src_data_431(\mm_interconnect_0|cmd_mux_001|src_data[43]~combout ),
	.src_data_421(\mm_interconnect_0|cmd_mux_001|src_data[42]~combout ),
	.src_data_401(\mm_interconnect_0|cmd_mux_001|src_data[40]~combout ),
	.src_data_391(\mm_interconnect_0|cmd_mux_001|src_data[39]~combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_001|src_payload~1_combout ),
	.src_data_321(\mm_interconnect_0|cmd_mux_001|src_data[32]~combout ),
	.av_readdata_8(\jtag_uart_0|av_readdata[8]~0_combout ),
	.d_writedata_27(\nios2_gen2_0|cpu|d_writedata[27]~q ),
	.src_payload31(\mm_interconnect_0|cmd_mux_002|src_payload~27_combout ),
	.d_writedata_28(\nios2_gen2_0|cpu|d_writedata[28]~q ),
	.src_payload32(\mm_interconnect_0|cmd_mux_002|src_payload~28_combout ),
	.d_writedata_29(\nios2_gen2_0|cpu|d_writedata[29]~q ),
	.src_payload33(\mm_interconnect_0|cmd_mux_002|src_payload~29_combout ),
	.d_writedata_30(\nios2_gen2_0|cpu|d_writedata[30]~q ),
	.src_payload34(\mm_interconnect_0|cmd_mux_002|src_payload~30_combout ),
	.d_writedata_31(\nios2_gen2_0|cpu|d_writedata[31]~q ),
	.src_payload35(\mm_interconnect_0|cmd_mux_002|src_payload~31_combout ),
	.ac(\jtag_uart_0|ac~q ),
	.av_readdata_9(\jtag_uart_0|av_readdata[9]~combout ),
	.b_full1(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.woverflow(\jtag_uart_0|woverflow~q ),
	.rvalid(\jtag_uart_0|rvalid~q ),
	.src_payload36(\mm_interconnect_0|rsp_mux|src_payload~2_combout ),
	.src_payload37(\mm_interconnect_0|cmd_mux_001|src_payload~2_combout ),
	.src_payload38(\mm_interconnect_0|rsp_mux|src_payload~3_combout ),
	.src_payload39(\mm_interconnect_0|rsp_mux|src_payload~4_combout ),
	.src_payload40(\mm_interconnect_0|rsp_mux|src_payload~5_combout ),
	.src_payload41(\mm_interconnect_0|rsp_mux|src_payload~6_combout ),
	.src_payload42(\mm_interconnect_0|rsp_mux|src_payload~7_combout ),
	.src_payload43(\mm_interconnect_0|rsp_mux|src_payload~8_combout ),
	.src_payload44(\mm_interconnect_0|rsp_mux|src_payload~9_combout ),
	.src_payload45(\mm_interconnect_0|cmd_mux_001|src_payload~3_combout ),
	.src_payload46(\mm_interconnect_0|cmd_mux_001|src_payload~4_combout ),
	.src_payload47(\mm_interconnect_0|cmd_mux_001|src_payload~5_combout ),
	.src_data_341(\mm_interconnect_0|cmd_mux_001|src_data[34]~combout ),
	.src_payload48(\mm_interconnect_0|cmd_mux_001|src_payload~6_combout ),
	.src_payload49(\mm_interconnect_0|cmd_mux_001|src_payload~7_combout ),
	.src_data_351(\mm_interconnect_0|cmd_mux_001|src_data[35]~combout ),
	.src_payload50(\mm_interconnect_0|cmd_mux_001|src_payload~8_combout ),
	.src_payload51(\mm_interconnect_0|cmd_mux_001|src_payload~9_combout ),
	.src_payload52(\mm_interconnect_0|cmd_mux_001|src_payload~10_combout ),
	.src_data_331(\mm_interconnect_0|cmd_mux_001|src_data[33]~combout ),
	.src_payload53(\mm_interconnect_0|cmd_mux_001|src_payload~11_combout ),
	.src_payload54(\mm_interconnect_0|cmd_mux_001|src_payload~12_combout ),
	.src_payload55(\mm_interconnect_0|cmd_mux_001|src_payload~13_combout ),
	.src_payload56(\mm_interconnect_0|cmd_mux_001|src_payload~14_combout ),
	.src_payload57(\mm_interconnect_0|cmd_mux_001|src_payload~15_combout ),
	.src_payload58(\mm_interconnect_0|cmd_mux_001|src_payload~16_combout ),
	.src_payload59(\mm_interconnect_0|cmd_mux_001|src_payload~17_combout ),
	.src_payload60(\mm_interconnect_0|cmd_mux_001|src_payload~18_combout ),
	.src_payload61(\mm_interconnect_0|cmd_mux_001|src_payload~19_combout ),
	.src_payload62(\mm_interconnect_0|cmd_mux_001|src_payload~20_combout ),
	.src_payload63(\mm_interconnect_0|cmd_mux_001|src_payload~21_combout ),
	.src_payload64(\mm_interconnect_0|cmd_mux_001|src_payload~22_combout ),
	.src_payload65(\mm_interconnect_0|cmd_mux_001|src_payload~23_combout ),
	.src_payload66(\mm_interconnect_0|cmd_mux_001|src_payload~24_combout ),
	.src_payload67(\mm_interconnect_0|cmd_mux_001|src_payload~25_combout ),
	.src_payload68(\mm_interconnect_0|cmd_mux_001|src_payload~26_combout ),
	.src_payload69(\mm_interconnect_0|cmd_mux_001|src_payload~27_combout ),
	.src_payload70(\mm_interconnect_0|cmd_mux_001|src_payload~28_combout ),
	.src_payload71(\mm_interconnect_0|cmd_mux_001|src_payload~29_combout ),
	.src_payload72(\mm_interconnect_0|cmd_mux_001|src_payload~30_combout ),
	.src_payload73(\mm_interconnect_0|cmd_mux_001|src_payload~31_combout ),
	.src_payload74(\mm_interconnect_0|cmd_mux_001|src_payload~32_combout ),
	.GND_port(\~GND~combout ),
	.clk_clk(\clk_clk~input_o ));

niosLab2_niosLab2_pio_0 pio_0(
	.W_alu_result_4(\nios2_gen2_0|cpu|W_alu_result[4]~q ),
	.W_alu_result_3(\nios2_gen2_0|cpu|W_alu_result[3]~q ),
	.W_alu_result_2(\nios2_gen2_0|cpu|W_alu_result[2]~q ),
	.data_out_0(\pio_0|data_out[0]~q ),
	.data_out_1(\pio_0|data_out[1]~q ),
	.data_out_2(\pio_0|data_out[2]~q ),
	.data_out_3(\pio_0|data_out[3]~q ),
	.data_out_4(\pio_0|data_out[4]~q ),
	.data_out_5(\pio_0|data_out[5]~q ),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\nios2_gen2_0|cpu|d_writedata[5]~q ,\nios2_gen2_0|cpu|d_writedata[4]~q ,\nios2_gen2_0|cpu|d_writedata[3]~q ,\nios2_gen2_0|cpu|d_writedata[2]~q ,\nios2_gen2_0|cpu|d_writedata[1]~q ,
\nios2_gen2_0|cpu|d_writedata[0]~q }),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.mem_used_1(\mm_interconnect_0|pio_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.Equal2(\mm_interconnect_0|router|Equal2~0_combout ),
	.Equal21(\mm_interconnect_0|router|Equal2~1_combout ),
	.rst1(\jtag_uart_0|niosLab2_jtag_uart_0_alt_jtag_atlantic|rst1~q ),
	.wait_latency_counter_1(\mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[0]~q ),
	.d_write(\nios2_gen2_0|cpu|d_write~q ),
	.write_accepted(\mm_interconnect_0|nios2_gen2_0_data_master_translator|write_accepted~q ),
	.always0(\pio_0|always0~3_combout ),
	.always01(\pio_0|always0~4_combout ),
	.readdata_0(\pio_0|readdata[0]~0_combout ),
	.readdata_1(\pio_0|readdata[1]~1_combout ),
	.readdata_2(\pio_0|readdata[2]~2_combout ),
	.readdata_3(\pio_0|readdata[3]~3_combout ),
	.readdata_4(\pio_0|readdata[4]~4_combout ),
	.readdata_5(\pio_0|readdata[5]~5_combout ),
	.clk(\clk_clk~input_o ));

niosLab2_niosLab2_onchip_memory2_0 onchip_memory2_0(
	.q_a_0(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_22(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_23(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_24(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_25(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_26(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_11(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_12(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_13(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_14(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_15(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_16(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_1(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_2(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_3(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_4(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_5(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_8(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_10(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_17(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_9(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_18(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_19(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_20(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_21(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_6(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_7(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_27(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_28(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_29(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_30(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_31(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[31] ),
	.always2(\jtag_uart_0|always2~0_combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ),
	.mem_used_1(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.src2_valid(\mm_interconnect_0|cmd_demux|src2_valid~0_combout ),
	.src_valid(\mm_interconnect_0|cmd_mux_002|src_valid~0_combout ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_002|src_payload~0_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_002|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_002|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_002|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_002|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_002|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_002|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_002|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_002|src_data[45]~combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_002|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_0|cmd_mux_002|src_data[47]~combout ),
	.src_data_48(\mm_interconnect_0|cmd_mux_002|src_data[48]~combout ),
	.src_data_49(\mm_interconnect_0|cmd_mux_002|src_data[49]~combout ),
	.src_data_50(\mm_interconnect_0|cmd_mux_002|src_data[50]~combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_002|src_data[32]~combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_002|src_payload~1_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_002|src_data[34]~combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_002|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_002|src_payload~3_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_002|src_data[35]~combout ),
	.src_payload4(\mm_interconnect_0|cmd_mux_002|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_002|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_002|src_payload~6_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_002|src_data[33]~combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_002|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_002|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_002|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_002|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_002|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_002|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_002|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_002|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_002|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_002|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_002|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_002|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_002|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_002|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_002|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_002|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_002|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_002|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_002|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_002|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_002|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_002|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_002|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_002|src_payload~30_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_002|src_payload~31_combout ),
	.clk_clk(\clk_clk~input_o ));

niosLab2_niosLab2_jtag_uart_0 jtag_uart_0(
	.W_alu_result_2(\nios2_gen2_0|cpu|W_alu_result[2]~q ),
	.q_b_0(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.d_writedata_10(\nios2_gen2_0|cpu|d_writedata[10]~q ),
	.q_b_1(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_7(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_6(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.Add1(\jtag_uart_0|Add1~1_sumout ),
	.Add11(\jtag_uart_0|Add1~5_sumout ),
	.Add12(\jtag_uart_0|Add1~9_sumout ),
	.Add13(\jtag_uart_0|Add1~13_sumout ),
	.Add14(\jtag_uart_0|Add1~17_sumout ),
	.Add15(\jtag_uart_0|Add1~21_sumout ),
	.Add16(\jtag_uart_0|Add1~25_sumout ),
	.adapted_tdo(\jtag_uart_0|niosLab2_jtag_uart_0_alt_jtag_atlantic|adapted_tdo~q ),
	.d_writedata_0(\nios2_gen2_0|cpu|d_writedata[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.Equal2(\mm_interconnect_0|router|Equal2~0_combout ),
	.Equal21(\mm_interconnect_0|router|Equal2~1_combout ),
	.rst1(\jtag_uart_0|niosLab2_jtag_uart_0_alt_jtag_atlantic|rst1~q ),
	.d_write(\nios2_gen2_0|cpu|d_write~q ),
	.write_accepted(\mm_interconnect_0|nios2_gen2_0_data_master_translator|write_accepted~q ),
	.d_writedata_1(\nios2_gen2_0|cpu|d_writedata[1]~q ),
	.d_writedata_2(\nios2_gen2_0|cpu|d_writedata[2]~q ),
	.d_writedata_3(\nios2_gen2_0|cpu|d_writedata[3]~q ),
	.d_writedata_4(\nios2_gen2_0|cpu|d_writedata[4]~q ),
	.d_writedata_5(\nios2_gen2_0|cpu|d_writedata[5]~q ),
	.d_read(\nios2_gen2_0|cpu|d_read~q ),
	.read_accepted(\mm_interconnect_0|nios2_gen2_0_data_master_translator|read_accepted~q ),
	.always2(\jtag_uart_0|always2~0_combout ),
	.Equal3(\mm_interconnect_0|router|Equal3~0_combout ),
	.mem_used_1(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest1(\jtag_uart_0|av_waitrequest~q ),
	.av_waitrequest2(\jtag_uart_0|av_waitrequest~0_combout ),
	.b_full(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.ien_AF1(\jtag_uart_0|ien_AF~q ),
	.read_01(\jtag_uart_0|read_0~q ),
	.d_writedata_6(\nios2_gen2_0|cpu|d_writedata[6]~q ),
	.d_writedata_7(\nios2_gen2_0|cpu|d_writedata[7]~q ),
	.ien_AE1(\jtag_uart_0|ien_AE~q ),
	.b_non_empty(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.counter_reg_bit_1(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_5(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.av_readdata_8(\jtag_uart_0|av_readdata[8]~0_combout ),
	.ac1(\jtag_uart_0|ac~q ),
	.av_readdata_9(\jtag_uart_0|av_readdata[9]~combout ),
	.b_full1(\jtag_uart_0|the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.woverflow1(\jtag_uart_0|woverflow~q ),
	.rvalid1(\jtag_uart_0|rvalid~q ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.splitter_nodes_receive_0_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.clr_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.irf_reg_0_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.clk_clk(\clk_clk~input_o ));

cyclonev_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~GND .extended_lut = "off";
defparam \~GND .lut_mask = 64'h0000000000000000;
defparam \~GND .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\altera_internal_jtag~TDIUTAP ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 64'hEDDEFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\altera_internal_jtag~TDIUTAP ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .lut_mask = 64'hFFFFB77BFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 .lut_mask = 64'hFFFBFFFFFFFEFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 .lut_mask = 64'hFFFFFFFF7FFFF7FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 .shared_arith = "off";

assign \clk_clk~input_o  = clk_clk;

assign \reset_reset_n~input_o  = reset_reset_n;

assign leds_export[0] = \pio_0|data_out[0]~q ;

assign leds_export[1] = \pio_0|data_out[1]~q ;

assign leds_export[2] = \pio_0|data_out[2]~q ;

assign leds_export[3] = \pio_0|data_out[3]~q ;

assign leds_export[4] = \pio_0|data_out[4]~q ;

assign leds_export[5] = \pio_0|data_out[5]~q ;

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

cyclonev_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 64'h6666666666666666;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 64'h9696969696969696;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 64'hFFFFFFEFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 (
	.dataa(!\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.dataf(!\altera_internal_jtag~TDIUTAP ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .lut_mask = 64'hEFFEFAFCEFFEFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(!\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|ir_out[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4 .lut_mask = 64'hF3FFFFFF77FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .lut_mask = 64'hFFFFFFACFFFFFFAC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .lut_mask = 64'hDF1FDF1FDF1FDF1F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 .lut_mask = 64'hFDF7FFFFF7FDFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3 .lut_mask = 64'hCF5FFFFFCF5FFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .lut_mask = 64'h6F9F9F6FFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 64'hF9FFF6FFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .lut_mask = 64'hFF7FFFDFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .lut_mask = 64'h7FFFF7FFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|ir_out[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .lut_mask = 64'hB77BFFFFB77BFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 64'hFFFFFFDFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .lut_mask = 64'h77DD77DD77DD77DD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .lut_mask = 64'hDD7777DDDD7777DD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .lut_mask = 64'h77DDDD77DD7777DD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .lut_mask = 64'hD77D7DD77DD7D77D;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .lut_mask = 64'hF6F9F9F6F6F9F9F6;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .lut_mask = 64'hDFFDFFFFDFFDFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .lut_mask = 64'hDEEDEDDEDEEDEDDE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(!\nios2_gen2_0|cpu|the_niosLab2_nios2_gen2_0_cpu_nios2_oci|the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[0]~q ),
	.datad(!\jtag_uart_0|niosLab2_jtag_uart_0_alt_jtag_atlantic|adapted_tdo~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .lut_mask = 64'hFFAAAAFFAAFFFFAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .lut_mask = 64'hFBFEFEFBFEFBFBFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .lut_mask = 64'hFFFFFEFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .lut_mask = 64'hAAFFFFAAAAFFFFAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .lut_mask = 64'hFFFFFEFFFFFFFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(!\altera_internal_jtag~TDIUTAP ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 64'hDF8FDF8FDF8FDF8F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .lut_mask = 64'hD8FFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .lut_mask = 64'hFFFFFFFFDF8FFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .lut_mask = 64'h6996699669966996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .lut_mask = 64'hF7B3FFFFF7B3FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .lut_mask = 64'hBFFFBF3FFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .lut_mask = 64'hFFFFFFFFFFFFFFBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .lut_mask = 64'hFFFFFFFFBFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

cyclonev_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|~GND .extended_lut = "off";
defparam \auto_hub|~GND .lut_mask = 64'h0000000000000000;
defparam \auto_hub|~GND .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .shared_arith = "off";

endmodule

module niosLab2_altera_reset_controller (
	r_sync_rst1,
	r_early_rst1,
	altera_reset_synchronizer_int_chain_1,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	r_sync_rst1;
output 	r_early_rst1;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[2]~q ;
wire \altera_reset_synchronizer_int_chain[3]~q ;
wire \altera_reset_synchronizer_int_chain[4]~0_combout ;
wire \altera_reset_synchronizer_int_chain[4]~q ;
wire \r_sync_rst_chain[3]~q ;
wire \r_sync_rst_chain~1_combout ;
wire \r_sync_rst_chain[2]~q ;
wire \r_sync_rst_chain~0_combout ;
wire \r_sync_rst_chain[1]~q ;
wire \WideOr0~0_combout ;
wire \always2~0_combout ;


niosLab2_altera_reset_synchronizer alt_rst_req_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.altera_reset_synchronizer_int_chain_1(altera_reset_synchronizer_int_chain_1),
	.clk(clk_clk));

niosLab2_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk(clk_clk),
	.reset_reset_n(reset_reset_n));

dffeas r_sync_rst(
	.clk(clk_clk),
	.d(\WideOr0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_sync_rst1),
	.prn(vcc));
defparam r_sync_rst.is_wysiwyg = "true";
defparam r_sync_rst.power_up = "low";

dffeas r_early_rst(
	.clk(clk_clk),
	.d(\always2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_early_rst1),
	.prn(vcc));
defparam r_early_rst.is_wysiwyg = "true";
defparam r_early_rst.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk_clk),
	.d(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[2] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[2]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[2] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[2] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[3]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[3] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[3] .power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[4]~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[4]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[4]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \altera_reset_synchronizer_int_chain[4]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[4] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[4]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[4] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[4] .power_up = "low";

dffeas \r_sync_rst_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[3]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[3] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[3] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~1 (
	.dataa(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datab(!\r_sync_rst_chain[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~1 .extended_lut = "off";
defparam \r_sync_rst_chain~1 .lut_mask = 64'h7777777777777777;
defparam \r_sync_rst_chain~1 .shared_arith = "off";

dffeas \r_sync_rst_chain[2] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[2]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[2] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[2] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datab(!\r_sync_rst_chain[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~0 .extended_lut = "off";
defparam \r_sync_rst_chain~0 .lut_mask = 64'h7777777777777777;
defparam \r_sync_rst_chain~0 .shared_arith = "off";

dffeas \r_sync_rst_chain[1] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[1]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[1] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[1] .power_up = "low";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!r_sync_rst1),
	.datab(!\altera_reset_synchronizer_int_chain[4]~q ),
	.datac(!\r_sync_rst_chain[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \always2~0 (
	.dataa(!\r_sync_rst_chain[2]~q ),
	.datab(!\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always2~0 .shared_arith = "off";

endmodule

module niosLab2_altera_reset_synchronizer (
	altera_reset_synchronizer_int_chain_out1,
	altera_reset_synchronizer_int_chain_1,
	clk)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(altera_reset_synchronizer_int_chain_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[1]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[1]~0 .lut_mask = 64'h0000000000000000;
defparam \altera_reset_synchronizer_int_chain[1]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(altera_reset_synchronizer_int_chain_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module niosLab2_altera_reset_synchronizer_1 (
	altera_reset_synchronizer_int_chain_out1,
	clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module niosLab2_niosLab2_jtag_uart_0 (
	W_alu_result_2,
	q_b_0,
	d_writedata_10,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_7,
	q_b_6,
	Add1,
	Add11,
	Add12,
	Add13,
	Add14,
	Add15,
	Add16,
	adapted_tdo,
	d_writedata_0,
	r_sync_rst,
	Equal2,
	Equal21,
	rst1,
	d_write,
	write_accepted,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_read,
	read_accepted,
	always2,
	Equal3,
	mem_used_1,
	av_waitrequest1,
	av_waitrequest2,
	b_full,
	ien_AF1,
	read_01,
	d_writedata_6,
	d_writedata_7,
	ien_AE1,
	b_non_empty,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	av_readdata_8,
	ac1,
	av_readdata_9,
	b_full1,
	woverflow1,
	rvalid1,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_2;
output 	q_b_0;
input 	d_writedata_10;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_7;
output 	q_b_6;
output 	Add1;
output 	Add11;
output 	Add12;
output 	Add13;
output 	Add14;
output 	Add15;
output 	Add16;
output 	adapted_tdo;
input 	d_writedata_0;
input 	r_sync_rst;
input 	Equal2;
input 	Equal21;
output 	rst1;
input 	d_write;
input 	write_accepted;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_read;
input 	read_accepted;
output 	always2;
input 	Equal3;
input 	mem_used_1;
output 	av_waitrequest1;
output 	av_waitrequest2;
output 	b_full;
output 	ien_AF1;
output 	read_01;
input 	d_writedata_6;
input 	d_writedata_7;
output 	ien_AE1;
output 	b_non_empty;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	av_readdata_8;
output 	ac1;
output 	av_readdata_9;
output 	b_full1;
output 	woverflow1;
output 	rvalid1;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \t_dav~q ;
wire \niosLab2_jtag_uart_0_alt_jtag_atlantic|rvalid0~q ;
wire \r_val~q ;
wire \niosLab2_jtag_uart_0_alt_jtag_atlantic|r_ena1~q ;
wire \fifo_wr~q ;
wire \the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \r_val~0_combout ;
wire \fifo_rd~1_combout ;
wire \niosLab2_jtag_uart_0_alt_jtag_atlantic|t_ena~reg0_q ;
wire \wr_rfifo~combout ;
wire \niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[0]~q ;
wire \niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[1]~q ;
wire \niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[2]~q ;
wire \niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[3]~q ;
wire \niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[4]~q ;
wire \niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[5]~q ;
wire \fifo_wr~0_combout ;
wire \the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \niosLab2_jtag_uart_0_alt_jtag_atlantic|t_pause~reg0_q ;
wire \niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[7]~q ;
wire \niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[6]~q ;
wire \Add1~2 ;
wire \Add1~6 ;
wire \Add1~10 ;
wire \Add1~14 ;
wire \Add1~18 ;
wire \Add1~22 ;
wire \av_waitrequest~1_combout ;
wire \av_waitrequest~2_combout ;
wire \av_waitrequest~3_combout ;
wire \always2~1_combout ;
wire \ien_AF~0_combout ;
wire \fifo_rd~0_combout ;
wire \fifo_rd~2_combout ;
wire \pause_irq~0_combout ;
wire \pause_irq~q ;
wire \Add0~22 ;
wire \Add0~26 ;
wire \Add0~18 ;
wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~17_sumout ;
wire \Add0~21_sumout ;
wire \Add0~25_sumout ;
wire \LessThan1~0_combout ;
wire \LessThan1~1_combout ;
wire \fifo_AF~q ;
wire \ac~0_combout ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \fifo_AE~q ;
wire \woverflow~0_combout ;
wire \rvalid~0_combout ;


niosLab2_niosLab2_jtag_uart_0_scfifo_r the_niosLab2_jtag_uart_0_scfifo_r(
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.r_sync_rst(r_sync_rst),
	.av_waitrequest(\av_waitrequest~1_combout ),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.fifo_rd(\fifo_rd~0_combout ),
	.fifo_rd1(\fifo_rd~1_combout ),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(\niosLab2_jtag_uart_0_alt_jtag_atlantic|t_ena~reg0_q ),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.wr_rfifo(\wr_rfifo~combout ),
	.wdata_0(\niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[0]~q ),
	.wdata_1(\niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[1]~q ),
	.wdata_2(\niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_3(\niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_4(\niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_5(\niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_7(\niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[7]~q ),
	.wdata_6(\niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[6]~q ),
	.clk_clk(clk_clk));

niosLab2_alt_jtag_atlantic niosLab2_jtag_uart_0_alt_jtag_atlantic(
	.r_dat({\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ,\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ,\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ,
\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ,\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ,\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ,
\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ,\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.adapted_tdo1(adapted_tdo),
	.rst_n(r_sync_rst),
	.rst11(rst1),
	.t_dav(\t_dav~q ),
	.rvalid01(\niosLab2_jtag_uart_0_alt_jtag_atlantic|rvalid0~q ),
	.r_val(\r_val~q ),
	.r_ena11(\niosLab2_jtag_uart_0_alt_jtag_atlantic|r_ena1~q ),
	.t_ena(\niosLab2_jtag_uart_0_alt_jtag_atlantic|t_ena~reg0_q ),
	.wdata_0(\niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[0]~q ),
	.wdata_1(\niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[1]~q ),
	.wdata_2(\niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_3(\niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_4(\niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_5(\niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[5]~q ),
	.t_pause(\niosLab2_jtag_uart_0_alt_jtag_atlantic|t_pause~reg0_q ),
	.wdata_7(\niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[7]~q ),
	.wdata_6(\niosLab2_jtag_uart_0_alt_jtag_atlantic|wdata[6]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.clr_reg(clr_reg),
	.state_3(state_3),
	.state_8(state_8),
	.irf_reg_0_1(irf_reg_0_1),
	.clk(clk_clk));

niosLab2_niosLab2_jtag_uart_0_scfifo_w the_niosLab2_jtag_uart_0_scfifo_w(
	.q_b_7(\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_0(\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.rvalid0(\niosLab2_jtag_uart_0_alt_jtag_atlantic|rvalid0~q ),
	.r_val(\r_val~q ),
	.r_ena1(\niosLab2_jtag_uart_0_alt_jtag_atlantic|r_ena1~q ),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.fifo_wr(\fifo_wr~q ),
	.b_non_empty(\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.r_val1(\r_val~0_combout ),
	.b_full(b_full1),
	.counter_reg_bit_0(\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_3(\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_5(\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.clk_clk(clk_clk));

dffeas t_dav(
	.clk(clk_clk),
	.d(b_full),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\t_dav~q ),
	.prn(vcc));
defparam t_dav.is_wysiwyg = "true";
defparam t_dav.power_up = "low";

dffeas r_val(
	.clk(clk_clk),
	.d(\r_val~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_val~q ),
	.prn(vcc));
defparam r_val.is_wysiwyg = "true";
defparam r_val.power_up = "low";

dffeas fifo_wr(
	.clk(clk_clk),
	.d(\fifo_wr~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_wr~q ),
	.prn(vcc));
defparam fifo_wr.is_wysiwyg = "true";
defparam fifo_wr.power_up = "low";

cyclonev_lcell_comb \r_val~0 (
	.dataa(!\niosLab2_jtag_uart_0_alt_jtag_atlantic|rvalid0~q ),
	.datab(!\r_val~q ),
	.datac(!\niosLab2_jtag_uart_0_alt_jtag_atlantic|r_ena1~q ),
	.datad(!\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_val~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_val~0 .extended_lut = "off";
defparam \r_val~0 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \r_val~0 .shared_arith = "off";

cyclonev_lcell_comb \fifo_rd~1 (
	.dataa(!Equal2),
	.datab(!Equal21),
	.datac(!Equal3),
	.datad(!\av_waitrequest~3_combout ),
	.datae(!b_non_empty),
	.dataf(!\fifo_rd~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_rd~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_rd~1 .extended_lut = "off";
defparam \fifo_rd~1 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \fifo_rd~1 .shared_arith = "off";

cyclonev_lcell_comb wr_rfifo(
	.dataa(!b_full),
	.datab(!\niosLab2_jtag_uart_0_alt_jtag_atlantic|t_ena~reg0_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_rfifo~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam wr_rfifo.extended_lut = "off";
defparam wr_rfifo.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam wr_rfifo.shared_arith = "off";

cyclonev_lcell_comb \fifo_wr~0 (
	.dataa(!W_alu_result_2),
	.datab(!\av_waitrequest~1_combout ),
	.datac(!\always2~1_combout ),
	.datad(!b_full1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr~0 .extended_lut = "off";
defparam \fifo_wr~0 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \fifo_wr~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Add1),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h000000000000FF00;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add11),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h000000000000FF00;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add12),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h000000000000FF00;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add13),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h000000000000FF00;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add14),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h000000000000FF00;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add15),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h000000000000FF00;
defparam \Add1~21 .shared_arith = "off";

cyclonev_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b_full1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add16),
	.cout(),
	.shareout());
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h000000000000FF00;
defparam \Add1~25 .shared_arith = "off";

cyclonev_lcell_comb \always2~0 (
	.dataa(!d_write),
	.datab(!write_accepted),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always2),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always2~0 .shared_arith = "off";

dffeas av_waitrequest(
	.clk(clk_clk),
	.d(\av_waitrequest~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_waitrequest1),
	.prn(vcc));
defparam av_waitrequest.is_wysiwyg = "true";
defparam av_waitrequest.power_up = "low";

cyclonev_lcell_comb \av_waitrequest~0 (
	.dataa(!rst1),
	.datab(!d_write),
	.datac(!write_accepted),
	.datad(!d_read),
	.datae(!read_accepted),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest2),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest~0 .extended_lut = "off";
defparam \av_waitrequest~0 .lut_mask = 64'hFFFFF7FFFFFFF7FF;
defparam \av_waitrequest~0 .shared_arith = "off";

dffeas ien_AF(
	.clk(clk_clk),
	.d(d_writedata_0),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AF~0_combout ),
	.q(ien_AF1),
	.prn(vcc));
defparam ien_AF.is_wysiwyg = "true";
defparam ien_AF.power_up = "low";

dffeas read_0(
	.clk(clk_clk),
	.d(\fifo_rd~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_01),
	.prn(vcc));
defparam read_0.is_wysiwyg = "true";
defparam read_0.power_up = "low";

dffeas ien_AE(
	.clk(clk_clk),
	.d(d_writedata_1),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AF~0_combout ),
	.q(ien_AE1),
	.prn(vcc));
defparam ien_AE.is_wysiwyg = "true";
defparam ien_AE.power_up = "low";

cyclonev_lcell_comb \av_readdata[8]~0 (
	.dataa(!ien_AF1),
	.datab(!\pause_irq~q ),
	.datac(!\fifo_AF~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_readdata_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdata[8]~0 .extended_lut = "off";
defparam \av_readdata[8]~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \av_readdata[8]~0 .shared_arith = "off";

dffeas ac(
	.clk(clk_clk),
	.d(\ac~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ac1),
	.prn(vcc));
defparam ac.is_wysiwyg = "true";
defparam ac.power_up = "low";

cyclonev_lcell_comb \av_readdata[9] (
	.dataa(!ien_AE1),
	.datab(!\fifo_AE~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_readdata_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdata[9] .extended_lut = "off";
defparam \av_readdata[9] .lut_mask = 64'h7777777777777777;
defparam \av_readdata[9] .shared_arith = "off";

dffeas woverflow(
	.clk(clk_clk),
	.d(\woverflow~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(woverflow1),
	.prn(vcc));
defparam woverflow.is_wysiwyg = "true";
defparam woverflow.power_up = "low";

dffeas rvalid(
	.clk(clk_clk),
	.d(\rvalid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rvalid1),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

cyclonev_lcell_comb \av_waitrequest~1 (
	.dataa(!Equal2),
	.datab(!Equal21),
	.datac(!Equal3),
	.datad(!mem_used_1),
	.datae(!av_waitrequest1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_waitrequest~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest~1 .extended_lut = "off";
defparam \av_waitrequest~1 .lut_mask = 64'hFFFFFF7FFFFFFF7F;
defparam \av_waitrequest~1 .shared_arith = "off";

cyclonev_lcell_comb \av_waitrequest~2 (
	.dataa(!av_waitrequest2),
	.datab(!\av_waitrequest~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_waitrequest~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest~2 .extended_lut = "off";
defparam \av_waitrequest~2 .lut_mask = 64'h7777777777777777;
defparam \av_waitrequest~2 .shared_arith = "off";

cyclonev_lcell_comb \av_waitrequest~3 (
	.dataa(!mem_used_1),
	.datab(!av_waitrequest1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_waitrequest~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest~3 .extended_lut = "off";
defparam \av_waitrequest~3 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \av_waitrequest~3 .shared_arith = "off";

cyclonev_lcell_comb \always2~1 (
	.dataa(!rst1),
	.datab(!d_write),
	.datac(!write_accepted),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~1 .extended_lut = "off";
defparam \always2~1 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \always2~1 .shared_arith = "off";

cyclonev_lcell_comb \ien_AF~0 (
	.dataa(!Equal2),
	.datab(!Equal21),
	.datac(!W_alu_result_2),
	.datad(!Equal3),
	.datae(!\av_waitrequest~3_combout ),
	.dataf(!\always2~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ien_AF~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ien_AF~0 .extended_lut = "off";
defparam \ien_AF~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \ien_AF~0 .shared_arith = "off";

cyclonev_lcell_comb \fifo_rd~0 (
	.dataa(!rst1),
	.datab(!W_alu_result_2),
	.datac(!d_read),
	.datad(!read_accepted),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_rd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_rd~0 .extended_lut = "off";
defparam \fifo_rd~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \fifo_rd~0 .shared_arith = "off";

cyclonev_lcell_comb \fifo_rd~2 (
	.dataa(!Equal2),
	.datab(!Equal21),
	.datac(!Equal3),
	.datad(!\av_waitrequest~3_combout ),
	.datae(!\fifo_rd~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_rd~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_rd~2 .extended_lut = "off";
defparam \fifo_rd~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \fifo_rd~2 .shared_arith = "off";

cyclonev_lcell_comb \pause_irq~0 (
	.dataa(!read_01),
	.datab(!b_non_empty),
	.datac(!\pause_irq~q ),
	.datad(!\niosLab2_jtag_uart_0_alt_jtag_atlantic|t_pause~reg0_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pause_irq~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pause_irq~0 .extended_lut = "off";
defparam \pause_irq~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \pause_irq~0 .shared_arith = "off";

dffeas pause_irq(
	.clk(clk_clk),
	.d(\pause_irq~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pause_irq~q ),
	.prn(vcc));
defparam pause_irq.is_wysiwyg = "true";
defparam pause_irq.power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(!counter_reg_bit_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000000000FF00;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000000000FF00;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000000000FF00;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b_full),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000000000FF00;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000000000000000;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \LessThan1~0 (
	.dataa(!counter_reg_bit_0),
	.datab(!\Add0~17_sumout ),
	.datac(!\Add0~21_sumout ),
	.datad(!\Add0~25_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~0 .extended_lut = "off";
defparam \LessThan1~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan1~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan1~1 (
	.dataa(!\Add0~1_sumout ),
	.datab(!\Add0~5_sumout ),
	.datac(!\Add0~9_sumout ),
	.datad(!\Add0~13_sumout ),
	.datae(!\LessThan1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~1 .extended_lut = "off";
defparam \LessThan1~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \LessThan1~1 .shared_arith = "off";

dffeas fifo_AF(
	.clk(clk_clk),
	.d(\LessThan1~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AF~q ),
	.prn(vcc));
defparam fifo_AF.is_wysiwyg = "true";
defparam fifo_AF.power_up = "low";

cyclonev_lcell_comb \ac~0 (
	.dataa(!d_writedata_10),
	.datab(!\niosLab2_jtag_uart_0_alt_jtag_atlantic|t_ena~reg0_q ),
	.datac(!\ien_AF~0_combout ),
	.datad(!ac1),
	.datae(!\niosLab2_jtag_uart_0_alt_jtag_atlantic|t_pause~reg0_q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac~0 .extended_lut = "off";
defparam \ac~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \ac~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.datab(!\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.datac(!\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.datad(!\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!b_full1),
	.datab(!\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.datac(!\the_niosLab2_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.datad(!\LessThan0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \LessThan0~1 .shared_arith = "off";

dffeas fifo_AE(
	.clk(clk_clk),
	.d(\LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AE~q ),
	.prn(vcc));
defparam fifo_AE.is_wysiwyg = "true";
defparam fifo_AE.power_up = "low";

cyclonev_lcell_comb \woverflow~0 (
	.dataa(!W_alu_result_2),
	.datab(!\av_waitrequest~1_combout ),
	.datac(!\always2~1_combout ),
	.datad(!b_full1),
	.datae(!woverflow1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\woverflow~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \woverflow~0 .extended_lut = "off";
defparam \woverflow~0 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \woverflow~0 .shared_arith = "off";

cyclonev_lcell_comb \rvalid~0 (
	.dataa(!b_non_empty),
	.datab(!\fifo_rd~2_combout ),
	.datac(!rvalid1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rvalid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rvalid~0 .extended_lut = "off";
defparam \rvalid~0 .lut_mask = 64'h4747474747474747;
defparam \rvalid~0 .shared_arith = "off";

endmodule

module niosLab2_alt_jtag_atlantic (
	r_dat,
	adapted_tdo1,
	rst_n,
	rst11,
	t_dav,
	rvalid01,
	r_val,
	r_ena11,
	t_ena,
	wdata_0,
	wdata_1,
	wdata_2,
	wdata_3,
	wdata_4,
	wdata_5,
	t_pause,
	wdata_7,
	wdata_6,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[7:0] r_dat;
output 	adapted_tdo1;
input 	rst_n;
output 	rst11;
input 	t_dav;
output 	rvalid01;
input 	r_val;
output 	r_ena11;
output 	t_ena;
output 	wdata_0;
output 	wdata_1;
output 	wdata_2;
output 	wdata_3;
output 	wdata_4;
output 	wdata_5;
output 	t_pause;
output 	wdata_7;
output 	wdata_6;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \state~1_combout ;
wire \state~q ;
wire \td_shift[0]~2_combout ;
wire \count[2]~q ;
wire \count[3]~q ;
wire \count[4]~q ;
wire \count[5]~q ;
wire \count[6]~q ;
wire \count[7]~q ;
wire \count[8]~q ;
wire \count[9]~0_combout ;
wire \count[9]~q ;
wire \count[9]~_wirecell_combout ;
wire \count[0]~q ;
wire \count[1]~q ;
wire \state~0_combout ;
wire \user_saw_rvalid~0_combout ;
wire \user_saw_rvalid~q ;
wire \td_shift[10]~q ;
wire \r_ena~0_combout ;
wire \rdata[7]~q ;
wire \td_shift~3_combout ;
wire \td_shift[9]~q ;
wire \td_shift~0_combout ;
wire \tck_t_dav~0_combout ;
wire \tck_t_dav~q ;
wire \write_stalled~0_combout ;
wire \write_stalled~1_combout ;
wire \write_stalled~q ;
wire \td_shift~4_combout ;
wire \rdata[0]~q ;
wire \rdata[6]~q ;
wire \td_shift~12_combout ;
wire \td_shift[8]~q ;
wire \rdata[5]~q ;
wire \td_shift~11_combout ;
wire \td_shift[7]~q ;
wire \rdata[4]~q ;
wire \td_shift~10_combout ;
wire \td_shift[6]~q ;
wire \rdata[3]~q ;
wire \td_shift~9_combout ;
wire \td_shift[5]~q ;
wire \rdata[2]~q ;
wire \td_shift~8_combout ;
wire \td_shift[4]~q ;
wire \rdata[1]~q ;
wire \td_shift~7_combout ;
wire \td_shift[3]~q ;
wire \td_shift~6_combout ;
wire \td_shift[2]~q ;
wire \td_shift~5_combout ;
wire \td_shift[1]~q ;
wire \rvalid~q ;
wire \td_shift~1_combout ;
wire \td_shift[0]~q ;
wire \rvalid0~0_combout ;
wire \read_req~q ;
wire \read~0_combout ;
wire \read~q ;
wire \read1~q ;
wire \read2~q ;
wire \rst2~q ;
wire \rvalid0~1_combout ;
wire \write~0_combout ;
wire \wdata[1]~0_combout ;
wire \write~q ;
wire \write1~q ;
wire \write2~q ;
wire \always2~0_combout ;
wire \write_valid~q ;
wire \t_ena~0_combout ;
wire \jupdate~0_combout ;
wire \jupdate~q ;
wire \jupdate1~q ;
wire \jupdate2~q ;
wire \always2~1_combout ;
wire \t_pause~0_combout ;


dffeas adapted_tdo(
	.clk(!altera_internal_jtag),
	.d(\td_shift[0]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(adapted_tdo1),
	.prn(vcc));
defparam adapted_tdo.is_wysiwyg = "true";
defparam adapted_tdo.power_up = "low";

dffeas rst1(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rst11),
	.prn(vcc));
defparam rst1.is_wysiwyg = "true";
defparam rst1.power_up = "low";

dffeas rvalid0(
	.clk(clk),
	.d(\rvalid0~1_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rvalid01),
	.prn(vcc));
defparam rvalid0.is_wysiwyg = "true";
defparam rvalid0.power_up = "low";

dffeas r_ena1(
	.clk(clk),
	.d(\rvalid0~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_ena11),
	.prn(vcc));
defparam r_ena1.is_wysiwyg = "true";
defparam r_ena1.power_up = "low";

dffeas \t_ena~reg0 (
	.clk(clk),
	.d(\t_ena~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_ena),
	.prn(vcc));
defparam \t_ena~reg0 .is_wysiwyg = "true";
defparam \t_ena~reg0 .power_up = "low";

dffeas \wdata[0] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(wdata_0),
	.prn(vcc));
defparam \wdata[0] .is_wysiwyg = "true";
defparam \wdata[0] .power_up = "low";

dffeas \wdata[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift[5]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~0_combout ),
	.q(wdata_1),
	.prn(vcc));
defparam \wdata[1] .is_wysiwyg = "true";
defparam \wdata[1] .power_up = "low";

dffeas \wdata[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift[6]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~0_combout ),
	.q(wdata_2),
	.prn(vcc));
defparam \wdata[2] .is_wysiwyg = "true";
defparam \wdata[2] .power_up = "low";

dffeas \wdata[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift[7]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~0_combout ),
	.q(wdata_3),
	.prn(vcc));
defparam \wdata[3] .is_wysiwyg = "true";
defparam \wdata[3] .power_up = "low";

dffeas \wdata[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift[8]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~0_combout ),
	.q(wdata_4),
	.prn(vcc));
defparam \wdata[4] .is_wysiwyg = "true";
defparam \wdata[4] .power_up = "low";

dffeas \wdata[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~0_combout ),
	.q(wdata_5),
	.prn(vcc));
defparam \wdata[5] .is_wysiwyg = "true";
defparam \wdata[5] .power_up = "low";

dffeas \t_pause~reg0 (
	.clk(clk),
	.d(\t_pause~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_pause),
	.prn(vcc));
defparam \t_pause~reg0 .is_wysiwyg = "true";
defparam \t_pause~reg0 .power_up = "low";

dffeas \wdata[7] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~0_combout ),
	.q(wdata_7),
	.prn(vcc));
defparam \wdata[7] .is_wysiwyg = "true";
defparam \wdata[7] .power_up = "low";

dffeas \wdata[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~0_combout ),
	.q(wdata_6),
	.prn(vcc));
defparam \wdata[6] .is_wysiwyg = "true";
defparam \wdata[6] .power_up = "low";

cyclonev_lcell_comb \state~1 (
	.dataa(!splitter_nodes_receive_0_3),
	.datab(!virtual_ir_scan_reg),
	.datac(!state_3),
	.datad(!state_4),
	.datae(!\state~q ),
	.dataf(!altera_internal_jtag1),
	.datag(!irf_reg_0_1),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~1 .extended_lut = "on";
defparam \state~1 .lut_mask = 64'hFF6FFF6FFF6FFF6F;
defparam \state~1 .shared_arith = "off";

dffeas state(
	.clk(altera_internal_jtag),
	.d(\state~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state~q ),
	.prn(vcc));
defparam state.is_wysiwyg = "true";
defparam state.power_up = "low";

cyclonev_lcell_comb \td_shift[0]~2 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_0_3),
	.datad(!state_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift[0]~2 .extended_lut = "off";
defparam \td_shift[0]~2 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \td_shift[0]~2 .shared_arith = "off";

dffeas \count[2] (
	.clk(altera_internal_jtag),
	.d(\count[1]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

dffeas \count[3] (
	.clk(altera_internal_jtag),
	.d(\count[2]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

dffeas \count[4] (
	.clk(altera_internal_jtag),
	.d(\count[3]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

dffeas \count[5] (
	.clk(altera_internal_jtag),
	.d(\count[4]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

dffeas \count[6] (
	.clk(altera_internal_jtag),
	.d(\count[5]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[6]~q ),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

dffeas \count[7] (
	.clk(altera_internal_jtag),
	.d(\count[6]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[7]~q ),
	.prn(vcc));
defparam \count[7] .is_wysiwyg = "true";
defparam \count[7] .power_up = "low";

dffeas \count[8] (
	.clk(altera_internal_jtag),
	.d(\count[7]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[8]~q ),
	.prn(vcc));
defparam \count[8] .is_wysiwyg = "true";
defparam \count[8] .power_up = "low";

cyclonev_lcell_comb \count[9]~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!altera_internal_jtag1),
	.datad(!state_4),
	.datae(!\count[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count[9]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count[9]~0 .extended_lut = "off";
defparam \count[9]~0 .lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam \count[9]~0 .shared_arith = "off";

dffeas \count[9] (
	.clk(altera_internal_jtag),
	.d(\count[9]~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[9]~q ),
	.prn(vcc));
defparam \count[9] .is_wysiwyg = "true";
defparam \count[9] .power_up = "low";

cyclonev_lcell_comb \count[9]~_wirecell (
	.dataa(!\count[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count[9]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count[9]~_wirecell .extended_lut = "off";
defparam \count[9]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \count[9]~_wirecell .shared_arith = "off";

dffeas \count[0] (
	.clk(altera_internal_jtag),
	.d(\count[9]~_wirecell_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

dffeas \count[1] (
	.clk(altera_internal_jtag),
	.d(\count[0]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cyclonev_lcell_comb \state~0 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_0_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~0 .extended_lut = "off";
defparam \state~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \state~0 .shared_arith = "off";

cyclonev_lcell_comb \user_saw_rvalid~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\td_shift[0]~q ),
	.datac(!\state~q ),
	.datad(!\user_saw_rvalid~q ),
	.datae(!\state~0_combout ),
	.dataf(!\count[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_saw_rvalid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_saw_rvalid~0 .extended_lut = "off";
defparam \user_saw_rvalid~0 .lut_mask = 64'h7BFFB7FFB7FF7BFF;
defparam \user_saw_rvalid~0 .shared_arith = "off";

dffeas user_saw_rvalid(
	.clk(altera_internal_jtag),
	.d(\user_saw_rvalid~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\user_saw_rvalid~q ),
	.prn(vcc));
defparam user_saw_rvalid.is_wysiwyg = "true";
defparam user_saw_rvalid.power_up = "low";

dffeas \td_shift[10] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[10]~q ),
	.prn(vcc));
defparam \td_shift[10] .is_wysiwyg = "true";
defparam \td_shift[10] .power_up = "low";

cyclonev_lcell_comb \r_ena~0 (
	.dataa(!r_val),
	.datab(!r_ena11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_ena~0 .extended_lut = "off";
defparam \r_ena~0 .lut_mask = 64'h7777777777777777;
defparam \r_ena~0 .shared_arith = "off";

dffeas \rdata[7] (
	.clk(clk),
	.d(r_dat[7]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[7]~q ),
	.prn(vcc));
defparam \rdata[7] .is_wysiwyg = "true";
defparam \rdata[7] .power_up = "low";

cyclonev_lcell_comb \td_shift~3 (
	.dataa(!\count[9]~q ),
	.datab(!\td_shift[10]~q ),
	.datac(!\rdata[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~3 .extended_lut = "off";
defparam \td_shift~3 .lut_mask = 64'h2727272727272727;
defparam \td_shift~3 .shared_arith = "off";

dffeas \td_shift[9] (
	.clk(altera_internal_jtag),
	.d(\td_shift~3_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[9]~q ),
	.prn(vcc));
defparam \td_shift[9] .is_wysiwyg = "true";
defparam \td_shift[9] .power_up = "low";

cyclonev_lcell_comb \td_shift~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!\count[1]~q ),
	.datad(!\user_saw_rvalid~q ),
	.datae(!\td_shift[9]~q ),
	.dataf(!altera_internal_jtag1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~0 .extended_lut = "off";
defparam \td_shift~0 .lut_mask = 64'hFFFFBF8FFFFFFFFF;
defparam \td_shift~0 .shared_arith = "off";

cyclonev_lcell_comb \tck_t_dav~0 (
	.dataa(!t_dav),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tck_t_dav~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tck_t_dav~0 .extended_lut = "off";
defparam \tck_t_dav~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \tck_t_dav~0 .shared_arith = "off";

dffeas tck_t_dav(
	.clk(altera_internal_jtag),
	.d(\tck_t_dav~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tck_t_dav~q ),
	.prn(vcc));
defparam tck_t_dav.is_wysiwyg = "true";
defparam tck_t_dav.power_up = "low";

cyclonev_lcell_comb \write_stalled~0 (
	.dataa(!altera_internal_jtag1),
	.datab(!\tck_t_dav~q ),
	.datac(!\td_shift[10]~q ),
	.datad(!\write_stalled~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_stalled~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_stalled~0 .extended_lut = "off";
defparam \write_stalled~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \write_stalled~0 .shared_arith = "off";

cyclonev_lcell_comb \write_stalled~1 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!\count[1]~q ),
	.datad(!state_4),
	.datae(!virtual_ir_scan_reg),
	.dataf(!splitter_nodes_receive_0_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_stalled~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_stalled~1 .extended_lut = "off";
defparam \write_stalled~1 .lut_mask = 64'hFFFFBFFFFFFFFFFF;
defparam \write_stalled~1 .shared_arith = "off";

dffeas write_stalled(
	.clk(altera_internal_jtag),
	.d(\write_stalled~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\write_stalled~q ),
	.prn(vcc));
defparam write_stalled.is_wysiwyg = "true";
defparam write_stalled.power_up = "low";

cyclonev_lcell_comb \td_shift~4 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!\count[1]~q ),
	.datad(!\user_saw_rvalid~q ),
	.datae(!\td_shift[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~4 .extended_lut = "off";
defparam \td_shift~4 .lut_mask = 64'hFFFFFFBFFFFFFFBF;
defparam \td_shift~4 .shared_arith = "off";

dffeas \rdata[0] (
	.clk(clk),
	.d(r_dat[0]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[0]~q ),
	.prn(vcc));
defparam \rdata[0] .is_wysiwyg = "true";
defparam \rdata[0] .power_up = "low";

dffeas \rdata[6] (
	.clk(clk),
	.d(r_dat[6]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[6]~q ),
	.prn(vcc));
defparam \rdata[6] .is_wysiwyg = "true";
defparam \rdata[6] .power_up = "low";

cyclonev_lcell_comb \td_shift~12 (
	.dataa(!\td_shift[9]~q ),
	.datab(!\count[9]~q ),
	.datac(!\rdata[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~12 .extended_lut = "off";
defparam \td_shift~12 .lut_mask = 64'h4747474747474747;
defparam \td_shift~12 .shared_arith = "off";

dffeas \td_shift[8] (
	.clk(altera_internal_jtag),
	.d(\td_shift~12_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[8]~q ),
	.prn(vcc));
defparam \td_shift[8] .is_wysiwyg = "true";
defparam \td_shift[8] .power_up = "low";

dffeas \rdata[5] (
	.clk(clk),
	.d(r_dat[5]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[5]~q ),
	.prn(vcc));
defparam \rdata[5] .is_wysiwyg = "true";
defparam \rdata[5] .power_up = "low";

cyclonev_lcell_comb \td_shift~11 (
	.dataa(!\count[9]~q ),
	.datab(!state_4),
	.datac(!\td_shift~4_combout ),
	.datad(!\td_shift[8]~q ),
	.datae(!\rdata[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~11 .extended_lut = "off";
defparam \td_shift~11 .lut_mask = 64'hB1FFFFFFB1FFFFFF;
defparam \td_shift~11 .shared_arith = "off";

dffeas \td_shift[7] (
	.clk(altera_internal_jtag),
	.d(\td_shift~11_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[7]~q ),
	.prn(vcc));
defparam \td_shift[7] .is_wysiwyg = "true";
defparam \td_shift[7] .power_up = "low";

dffeas \rdata[4] (
	.clk(clk),
	.d(r_dat[4]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[4]~q ),
	.prn(vcc));
defparam \rdata[4] .is_wysiwyg = "true";
defparam \rdata[4] .power_up = "low";

cyclonev_lcell_comb \td_shift~10 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\td_shift~4_combout ),
	.datae(!\td_shift[7]~q ),
	.dataf(!\rdata[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~10 .extended_lut = "off";
defparam \td_shift~10 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \td_shift~10 .shared_arith = "off";

dffeas \td_shift[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift~10_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[6]~q ),
	.prn(vcc));
defparam \td_shift[6] .is_wysiwyg = "true";
defparam \td_shift[6] .power_up = "low";

dffeas \rdata[3] (
	.clk(clk),
	.d(r_dat[3]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[3]~q ),
	.prn(vcc));
defparam \rdata[3] .is_wysiwyg = "true";
defparam \rdata[3] .power_up = "low";

cyclonev_lcell_comb \td_shift~9 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\td_shift~4_combout ),
	.datae(!\td_shift[6]~q ),
	.dataf(!\rdata[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~9 .extended_lut = "off";
defparam \td_shift~9 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \td_shift~9 .shared_arith = "off";

dffeas \td_shift[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift~9_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[5]~q ),
	.prn(vcc));
defparam \td_shift[5] .is_wysiwyg = "true";
defparam \td_shift[5] .power_up = "low";

dffeas \rdata[2] (
	.clk(clk),
	.d(r_dat[2]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[2]~q ),
	.prn(vcc));
defparam \rdata[2] .is_wysiwyg = "true";
defparam \rdata[2] .power_up = "low";

cyclonev_lcell_comb \td_shift~8 (
	.dataa(!\count[9]~q ),
	.datab(!state_4),
	.datac(!\td_shift~4_combout ),
	.datad(!\td_shift[5]~q ),
	.datae(!\rdata[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~8 .extended_lut = "off";
defparam \td_shift~8 .lut_mask = 64'hB1FFFFFFB1FFFFFF;
defparam \td_shift~8 .shared_arith = "off";

dffeas \td_shift[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift~8_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[4]~q ),
	.prn(vcc));
defparam \td_shift[4] .is_wysiwyg = "true";
defparam \td_shift[4] .power_up = "low";

dffeas \rdata[1] (
	.clk(clk),
	.d(r_dat[1]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[1]~q ),
	.prn(vcc));
defparam \rdata[1] .is_wysiwyg = "true";
defparam \rdata[1] .power_up = "low";

cyclonev_lcell_comb \td_shift~7 (
	.dataa(!\count[9]~q ),
	.datab(!state_4),
	.datac(!\td_shift~4_combout ),
	.datad(!\td_shift[4]~q ),
	.datae(!\rdata[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~7 .extended_lut = "off";
defparam \td_shift~7 .lut_mask = 64'hB1FFFFFFB1FFFFFF;
defparam \td_shift~7 .shared_arith = "off";

dffeas \td_shift[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift~7_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[3]~q ),
	.prn(vcc));
defparam \td_shift[3] .is_wysiwyg = "true";
defparam \td_shift[3] .power_up = "low";

cyclonev_lcell_comb \td_shift~6 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\td_shift~4_combout ),
	.datae(!\rdata[0]~q ),
	.dataf(!\td_shift[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~6 .extended_lut = "off";
defparam \td_shift~6 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \td_shift~6 .shared_arith = "off";

dffeas \td_shift[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift~6_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[2]~q ),
	.prn(vcc));
defparam \td_shift[2] .is_wysiwyg = "true";
defparam \td_shift[2] .power_up = "low";

cyclonev_lcell_comb \td_shift~5 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\write_stalled~q ),
	.datae(!\td_shift~4_combout ),
	.dataf(!\td_shift[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~5 .extended_lut = "off";
defparam \td_shift~5 .lut_mask = 64'hFFFF7DFFFFFFFFFF;
defparam \td_shift~5 .shared_arith = "off";

dffeas \td_shift[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift~5_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[1]~q ),
	.prn(vcc));
defparam \td_shift[1] .is_wysiwyg = "true";
defparam \td_shift[1] .power_up = "low";

dffeas rvalid(
	.clk(clk),
	.d(rvalid01),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rvalid~q ),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

cyclonev_lcell_comb \td_shift~1 (
	.dataa(!\state~q ),
	.datab(!\td_shift~0_combout ),
	.datac(!\tck_t_dav~q ),
	.datad(!\td_shift[1]~q ),
	.datae(!\count[9]~q ),
	.dataf(!\rvalid~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~1 .extended_lut = "off";
defparam \td_shift~1 .lut_mask = 64'hBFFFEFFFFFFFFFFF;
defparam \td_shift~1 .shared_arith = "off";

dffeas \td_shift[0] (
	.clk(altera_internal_jtag),
	.d(\td_shift~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[0]~q ),
	.prn(vcc));
defparam \td_shift[0] .is_wysiwyg = "true";
defparam \td_shift[0] .power_up = "low";

cyclonev_lcell_comb \rvalid0~0 (
	.dataa(!rvalid01),
	.datab(!r_val),
	.datac(!r_ena11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rvalid0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rvalid0~0 .extended_lut = "off";
defparam \rvalid0~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \rvalid0~0 .shared_arith = "off";

dffeas read_req(
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\read_req~q ),
	.prn(vcc));
defparam read_req.is_wysiwyg = "true";
defparam read_req.power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!\read~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \read~0 .shared_arith = "off";

dffeas read(
	.clk(altera_internal_jtag),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

dffeas read1(
	.clk(clk),
	.d(\read~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read1~q ),
	.prn(vcc));
defparam read1.is_wysiwyg = "true";
defparam read1.power_up = "low";

dffeas read2(
	.clk(clk),
	.d(\read1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read2~q ),
	.prn(vcc));
defparam read2.is_wysiwyg = "true";
defparam read2.power_up = "low";

dffeas rst2(
	.clk(clk),
	.d(rst11),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rst2~q ),
	.prn(vcc));
defparam rst2.is_wysiwyg = "true";
defparam rst2.power_up = "low";

cyclonev_lcell_comb \rvalid0~1 (
	.dataa(!\user_saw_rvalid~q ),
	.datab(!\rvalid0~0_combout ),
	.datac(!\read_req~q ),
	.datad(!\read1~q ),
	.datae(!\read2~q ),
	.dataf(!\rst2~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rvalid0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rvalid0~1 .extended_lut = "off";
defparam \rvalid0~1 .lut_mask = 64'hFFFFFFFFFEFFFFFE;
defparam \rvalid0~1 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!\write~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \wdata[1]~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!state_4),
	.datad(!virtual_ir_scan_reg),
	.datae(!splitter_nodes_receive_0_3),
	.dataf(!\count[8]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wdata[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wdata[1]~0 .extended_lut = "off";
defparam \wdata[1]~0 .lut_mask = 64'hFFBFFFFFFFFFFFFF;
defparam \wdata[1]~0 .shared_arith = "off";

dffeas write(
	.clk(altera_internal_jtag),
	.d(\write~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~0_combout ),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas write1(
	.clk(clk),
	.d(\write~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write1~q ),
	.prn(vcc));
defparam write1.is_wysiwyg = "true";
defparam write1.power_up = "low";

dffeas write2(
	.clk(clk),
	.d(\write1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write2~q ),
	.prn(vcc));
defparam write2.is_wysiwyg = "true";
defparam write2.power_up = "low";

cyclonev_lcell_comb \always2~0 (
	.dataa(!\write1~q ),
	.datab(!\write2~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'h6666666666666666;
defparam \always2~0 .shared_arith = "off";

dffeas write_valid(
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\write_valid~q ),
	.prn(vcc));
defparam write_valid.is_wysiwyg = "true";
defparam write_valid.power_up = "low";

cyclonev_lcell_comb \t_ena~0 (
	.dataa(!t_dav),
	.datab(!\write_stalled~q ),
	.datac(!\rst2~q ),
	.datad(!t_ena),
	.datae(!\always2~0_combout ),
	.dataf(!\write_valid~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\t_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \t_ena~0 .extended_lut = "off";
defparam \t_ena~0 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \t_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \jupdate~0 (
	.dataa(!irf_reg_0_1),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_0_3),
	.datad(!\jupdate~q ),
	.datae(!state_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jupdate~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jupdate~0 .extended_lut = "off";
defparam \jupdate~0 .lut_mask = 64'h9669699696696996;
defparam \jupdate~0 .shared_arith = "off";

dffeas jupdate(
	.clk(!altera_internal_jtag),
	.d(\jupdate~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate~q ),
	.prn(vcc));
defparam jupdate.is_wysiwyg = "true";
defparam jupdate.power_up = "low";

dffeas jupdate1(
	.clk(clk),
	.d(\jupdate~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate1~q ),
	.prn(vcc));
defparam jupdate1.is_wysiwyg = "true";
defparam jupdate1.power_up = "low";

dffeas jupdate2(
	.clk(clk),
	.d(\jupdate1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate2~q ),
	.prn(vcc));
defparam jupdate2.is_wysiwyg = "true";
defparam jupdate2.power_up = "low";

cyclonev_lcell_comb \always2~1 (
	.dataa(!\jupdate1~q ),
	.datab(!\jupdate2~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~1 .extended_lut = "off";
defparam \always2~1 .lut_mask = 64'h6666666666666666;
defparam \always2~1 .shared_arith = "off";

cyclonev_lcell_comb \t_pause~0 (
	.dataa(!t_dav),
	.datab(!\write_stalled~q ),
	.datac(!\rst2~q ),
	.datad(!\always2~0_combout ),
	.datae(!\write_valid~q ),
	.dataf(!\always2~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\t_pause~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \t_pause~0 .extended_lut = "off";
defparam \t_pause~0 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \t_pause~0 .shared_arith = "off";

endmodule

module niosLab2_niosLab2_jtag_uart_0_scfifo_r (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_7,
	q_b_6,
	r_sync_rst,
	av_waitrequest,
	b_full,
	b_non_empty,
	fifo_rd,
	fifo_rd1,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	wr_rfifo,
	wdata_0,
	wdata_1,
	wdata_2,
	wdata_3,
	wdata_4,
	wdata_5,
	wdata_7,
	wdata_6,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_7;
output 	q_b_6;
input 	r_sync_rst;
input 	av_waitrequest;
output 	b_full;
output 	b_non_empty;
input 	fifo_rd;
input 	fifo_rd1;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	wr_rfifo;
input 	wdata_0;
input 	wdata_1;
input 	wdata_2;
input 	wdata_3;
input 	wdata_4;
input 	wdata_5;
input 	wdata_7;
input 	wdata_6;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosLab2_scfifo_1 rfifo(
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.r_sync_rst(r_sync_rst),
	.av_waitrequest(av_waitrequest),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.fifo_rd(fifo_rd),
	.fifo_rd1(fifo_rd1),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.wrreq(wr_rfifo),
	.data({wdata_7,wdata_6,wdata_5,wdata_4,wdata_3,wdata_2,wdata_1,wdata_0}),
	.clock(clk_clk));

endmodule

module niosLab2_scfifo_1 (
	q,
	r_sync_rst,
	av_waitrequest,
	b_full,
	b_non_empty,
	fifo_rd,
	fifo_rd1,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	wrreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
input 	av_waitrequest;
output 	b_full;
output 	b_non_empty;
input 	fifo_rd;
input 	fifo_rd1;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	wrreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosLab2_scfifo_3291 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.r_sync_rst(r_sync_rst),
	.av_waitrequest(av_waitrequest),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.fifo_rd(fifo_rd),
	.fifo_rd1(fifo_rd1),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.wrreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock));

endmodule

module niosLab2_scfifo_3291 (
	q,
	r_sync_rst,
	av_waitrequest,
	b_full,
	b_non_empty,
	fifo_rd,
	fifo_rd1,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	wrreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
input 	av_waitrequest;
output 	b_full;
output 	b_non_empty;
input 	fifo_rd;
input 	fifo_rd1;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	wrreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosLab2_a_dpfifo_5771 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.r_sync_rst(r_sync_rst),
	.av_waitrequest(av_waitrequest),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.fifo_rd(fifo_rd),
	.fifo_rd1(fifo_rd1),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.wreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock));

endmodule

module niosLab2_a_dpfifo_5771 (
	q,
	r_sync_rst,
	av_waitrequest,
	b_full,
	b_non_empty,
	fifo_rd,
	fifo_rd1,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	wreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
input 	av_waitrequest;
output 	b_full;
output 	b_non_empty;
input 	fifo_rd;
input 	fifo_rd1;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	wreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


niosLab2_altsyncram_7pu1 FIFOram(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.clocken1(fifo_rd1),
	.wren_a(wreq),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.clock0(clock),
	.clock1(clock));

niosLab2_a_fefifo_7cf fifo_state(
	.r_sync_rst(r_sync_rst),
	.av_waitrequest(av_waitrequest),
	.b_full1(b_full),
	.b_non_empty1(b_non_empty),
	.fifo_rd(fifo_rd),
	.fifo_rd1(fifo_rd1),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.wr_rfifo(wreq),
	.clock(clock));

niosLab2_cntr_jgb_1 wr_ptr(
	.r_sync_rst(r_sync_rst),
	.wr_rfifo(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

niosLab2_cntr_jgb rd_ptr_count(
	.r_sync_rst(r_sync_rst),
	.fifo_rd(fifo_rd1),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

endmodule

module niosLab2_a_fefifo_7cf (
	r_sync_rst,
	av_waitrequest,
	b_full1,
	b_non_empty1,
	fifo_rd,
	fifo_rd1,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	wr_rfifo,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	av_waitrequest;
output 	b_full1;
output 	b_non_empty1;
input 	fifo_rd;
input 	fifo_rd1;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	wr_rfifo;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~2_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \b_non_empty~0_combout ;


niosLab2_cntr_vg7 count_usedw(
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.wr_rfifo(wr_rfifo),
	._(\_~2_combout ),
	.clock(clock));

cyclonev_lcell_comb \_~2 (
	.dataa(!av_waitrequest),
	.datab(!b_non_empty1),
	.datac(!fifo_rd),
	.datad(!wr_rfifo),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~2 .extended_lut = "off";
defparam \_~2 .lut_mask = 64'h6996699669966996;
defparam \_~2 .shared_arith = "off";

dffeas b_full(
	.clk(clock),
	.d(\b_full~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

cyclonev_lcell_comb \b_full~0 (
	.dataa(!b_non_empty1),
	.datab(!counter_reg_bit_5),
	.datac(!counter_reg_bit_4),
	.datad(!counter_reg_bit_3),
	.datae(!counter_reg_bit_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~0 .extended_lut = "off";
defparam \b_full~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \b_full~0 .shared_arith = "off";

cyclonev_lcell_comb \b_full~1 (
	.dataa(!b_full1),
	.datab(!fifo_rd1),
	.datac(!counter_reg_bit_1),
	.datad(!counter_reg_bit_0),
	.datae(!t_ena),
	.dataf(!\b_full~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~1 .extended_lut = "off";
defparam \b_full~1 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \b_full~1 .shared_arith = "off";

cyclonev_lcell_comb \_~0 (
	.dataa(!b_full1),
	.datab(!counter_reg_bit_5),
	.datac(!counter_reg_bit_4),
	.datad(!t_ena),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \_~0 .shared_arith = "off";

cyclonev_lcell_comb \_~1 (
	.dataa(!counter_reg_bit_3),
	.datab(!counter_reg_bit_2),
	.datac(!counter_reg_bit_1),
	.datad(!counter_reg_bit_0),
	.datae(!\_~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~1 .extended_lut = "off";
defparam \_~1 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \_~1 .shared_arith = "off";

cyclonev_lcell_comb \b_non_empty~0 (
	.dataa(!b_full1),
	.datab(!b_non_empty1),
	.datac(!fifo_rd1),
	.datad(!t_ena),
	.datae(!\_~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~0 .extended_lut = "off";
defparam \b_non_empty~0 .lut_mask = 64'hF7FFD5FFF7FFD5FF;
defparam \b_non_empty~0 .shared_arith = "off";

endmodule

module niosLab2_cntr_vg7 (
	r_sync_rst,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	wr_rfifo,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	wr_rfifo;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita2~sumout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module niosLab2_altsyncram_7pu1 (
	q_b,
	clocken1,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	clocken1;
input 	wren_a;
input 	[7:0] data_a;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "niosLab2_jtag_uart_0:jtag_uart_0|niosLab2_jtag_uart_0_scfifo_r:the_niosLab2_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "niosLab2_jtag_uart_0:jtag_uart_0|niosLab2_jtag_uart_0_scfifo_r:the_niosLab2_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "niosLab2_jtag_uart_0:jtag_uart_0|niosLab2_jtag_uart_0_scfifo_r:the_niosLab2_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "niosLab2_jtag_uart_0:jtag_uart_0|niosLab2_jtag_uart_0_scfifo_r:the_niosLab2_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "niosLab2_jtag_uart_0:jtag_uart_0|niosLab2_jtag_uart_0_scfifo_r:the_niosLab2_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "niosLab2_jtag_uart_0:jtag_uart_0|niosLab2_jtag_uart_0_scfifo_r:the_niosLab2_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "niosLab2_jtag_uart_0:jtag_uart_0|niosLab2_jtag_uart_0_scfifo_r:the_niosLab2_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "niosLab2_jtag_uart_0:jtag_uart_0|niosLab2_jtag_uart_0_scfifo_r:the_niosLab2_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

endmodule

module niosLab2_cntr_jgb (
	r_sync_rst,
	fifo_rd,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_rd;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module niosLab2_cntr_jgb_1 (
	r_sync_rst,
	wr_rfifo,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	wr_rfifo;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module niosLab2_niosLab2_jtag_uart_0_scfifo_w (
	q_b_7,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	d_writedata_0,
	r_sync_rst,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	rvalid0,
	r_val,
	r_ena1,
	d_writedata_6,
	d_writedata_7,
	fifo_wr,
	b_non_empty,
	r_val1,
	b_full,
	counter_reg_bit_0,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_7;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
input 	d_writedata_0;
input 	r_sync_rst;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	rvalid0;
input 	r_val;
input 	r_ena1;
input 	d_writedata_6;
input 	d_writedata_7;
input 	fifo_wr;
output 	b_non_empty;
input 	r_val1;
output 	b_full;
output 	counter_reg_bit_0;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosLab2_scfifo_2 wfifo(
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data({d_writedata_7,d_writedata_6,d_writedata_5,d_writedata_4,d_writedata_3,d_writedata_2,d_writedata_1,d_writedata_0}),
	.r_sync_rst(r_sync_rst),
	.rvalid0(rvalid0),
	.r_val(r_val),
	.r_ena1(r_ena1),
	.wrreq(fifo_wr),
	.b_non_empty(b_non_empty),
	.r_val1(r_val1),
	.b_full(b_full),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.clock(clk_clk));

endmodule

module niosLab2_scfifo_2 (
	q,
	data,
	r_sync_rst,
	rvalid0,
	r_val,
	r_ena1,
	wrreq,
	b_non_empty,
	r_val1,
	b_full,
	counter_reg_bit_0,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
input 	rvalid0;
input 	r_val;
input 	r_ena1;
input 	wrreq;
output 	b_non_empty;
input 	r_val1;
output 	b_full;
output 	counter_reg_bit_0;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosLab2_scfifo_3291_1 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.r_sync_rst(r_sync_rst),
	.rvalid0(rvalid0),
	.r_val(r_val),
	.r_ena1(r_ena1),
	.wrreq(wrreq),
	.b_non_empty(b_non_empty),
	.r_val1(r_val1),
	.b_full(b_full),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.clock(clock));

endmodule

module niosLab2_scfifo_3291_1 (
	q,
	data,
	r_sync_rst,
	rvalid0,
	r_val,
	r_ena1,
	wrreq,
	b_non_empty,
	r_val1,
	b_full,
	counter_reg_bit_0,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
input 	rvalid0;
input 	r_val;
input 	r_ena1;
input 	wrreq;
output 	b_non_empty;
input 	r_val1;
output 	b_full;
output 	counter_reg_bit_0;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosLab2_a_dpfifo_5771_1 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.r_sync_rst(r_sync_rst),
	.rvalid0(rvalid0),
	.r_val(r_val),
	.r_ena1(r_ena1),
	.wreq(wrreq),
	.b_non_empty(b_non_empty),
	.r_val1(r_val1),
	.b_full(b_full),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.clock(clock));

endmodule

module niosLab2_a_dpfifo_5771_1 (
	q,
	data,
	r_sync_rst,
	rvalid0,
	r_val,
	r_ena1,
	wreq,
	b_non_empty,
	r_val1,
	b_full,
	counter_reg_bit_0,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
input 	rvalid0;
input 	r_val;
input 	r_ena1;
input 	wreq;
output 	b_non_empty;
input 	r_val1;
output 	b_full;
output 	counter_reg_bit_0;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


niosLab2_cntr_jgb_3 wr_ptr(
	.r_sync_rst(r_sync_rst),
	.fifo_wr(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

niosLab2_cntr_jgb_2 rd_ptr_count(
	.r_sync_rst(r_sync_rst),
	.r_val(r_val1),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

niosLab2_altsyncram_7pu1_1 FIFOram(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.wren_a(wreq),
	.clocken1(r_val1),
	.address_a({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.clock0(clock),
	.clock1(clock));

niosLab2_a_fefifo_7cf_1 fifo_state(
	.r_sync_rst(r_sync_rst),
	.rvalid0(rvalid0),
	.r_val(r_val),
	.r_ena1(r_ena1),
	.fifo_wr(wreq),
	.b_non_empty1(b_non_empty),
	.r_val1(r_val1),
	.b_full1(b_full),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.clock(clock));

endmodule

module niosLab2_a_fefifo_7cf_1 (
	r_sync_rst,
	rvalid0,
	r_val,
	r_ena1,
	fifo_wr,
	b_non_empty1,
	r_val1,
	b_full1,
	counter_reg_bit_0,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	rvalid0;
input 	r_val;
input 	r_ena1;
input 	fifo_wr;
output 	b_non_empty1;
input 	r_val1;
output 	b_full1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~0_combout ;
wire \b_non_empty~0_combout ;
wire \b_non_empty~1_combout ;
wire \b_non_empty~2_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;


niosLab2_cntr_vg7_1 count_usedw(
	.r_sync_rst(r_sync_rst),
	.fifo_wr(fifo_wr),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	._(\_~0_combout ),
	.clock(clock));

cyclonev_lcell_comb \_~0 (
	.dataa(!rvalid0),
	.datab(!r_val),
	.datac(!r_ena1),
	.datad(!fifo_wr),
	.datae(!b_non_empty1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'h9669699696696996;
defparam \_~0 .shared_arith = "off";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

dffeas b_full(
	.clk(clock),
	.d(\b_full~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

cyclonev_lcell_comb \b_non_empty~0 (
	.dataa(!counter_reg_bit_2),
	.datab(!counter_reg_bit_1),
	.datac(!counter_reg_bit_5),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~0 .extended_lut = "off";
defparam \b_non_empty~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \b_non_empty~0 .shared_arith = "off";

cyclonev_lcell_comb \b_non_empty~1 (
	.dataa(!r_val1),
	.datab(!counter_reg_bit_0),
	.datac(!counter_reg_bit_3),
	.datad(!\b_non_empty~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~1 .extended_lut = "off";
defparam \b_non_empty~1 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \b_non_empty~1 .shared_arith = "off";

cyclonev_lcell_comb \b_non_empty~2 (
	.dataa(!fifo_wr),
	.datab(!b_non_empty1),
	.datac(!b_full1),
	.datad(!\b_non_empty~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~2 .extended_lut = "off";
defparam \b_non_empty~2 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \b_non_empty~2 .shared_arith = "off";

cyclonev_lcell_comb \b_full~0 (
	.dataa(!fifo_wr),
	.datab(!b_non_empty1),
	.datac(!counter_reg_bit_3),
	.datad(!counter_reg_bit_5),
	.datae(!counter_reg_bit_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~0 .extended_lut = "off";
defparam \b_full~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \b_full~0 .shared_arith = "off";

cyclonev_lcell_comb \b_full~1 (
	.dataa(!r_val1),
	.datab(!b_full1),
	.datac(!counter_reg_bit_0),
	.datad(!counter_reg_bit_2),
	.datae(!counter_reg_bit_1),
	.dataf(!\b_full~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~1 .extended_lut = "off";
defparam \b_full~1 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \b_full~1 .shared_arith = "off";

endmodule

module niosLab2_cntr_vg7_1 (
	r_sync_rst,
	fifo_wr,
	counter_reg_bit_0,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_wr;
output 	counter_reg_bit_0;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;
wire \counter_comb_bita4~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module niosLab2_altsyncram_7pu1_1 (
	q_b,
	data_a,
	wren_a,
	clocken1,
	address_a,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	[7:0] data_a;
input 	wren_a;
input 	clocken1;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "niosLab2_jtag_uart_0:jtag_uart_0|niosLab2_jtag_uart_0_scfifo_w:the_niosLab2_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "niosLab2_jtag_uart_0:jtag_uart_0|niosLab2_jtag_uart_0_scfifo_w:the_niosLab2_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "niosLab2_jtag_uart_0:jtag_uart_0|niosLab2_jtag_uart_0_scfifo_w:the_niosLab2_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "niosLab2_jtag_uart_0:jtag_uart_0|niosLab2_jtag_uart_0_scfifo_w:the_niosLab2_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "niosLab2_jtag_uart_0:jtag_uart_0|niosLab2_jtag_uart_0_scfifo_w:the_niosLab2_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "niosLab2_jtag_uart_0:jtag_uart_0|niosLab2_jtag_uart_0_scfifo_w:the_niosLab2_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "niosLab2_jtag_uart_0:jtag_uart_0|niosLab2_jtag_uart_0_scfifo_w:the_niosLab2_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "niosLab2_jtag_uart_0:jtag_uart_0|niosLab2_jtag_uart_0_scfifo_w:the_niosLab2_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

endmodule

module niosLab2_cntr_jgb_2 (
	r_sync_rst,
	r_val,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	r_val;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module niosLab2_cntr_jgb_3 (
	r_sync_rst,
	fifo_wr,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_wr;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module niosLab2_niosLab2_mm_interconnect_0 (
	W_alu_result_4,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_7,
	W_alu_result_6,
	W_alu_result_5,
	W_alu_result_12,
	W_alu_result_13,
	W_alu_result_14,
	W_alu_result_15,
	W_alu_result_16,
	W_alu_result_3,
	W_alu_result_2,
	F_pc_9,
	F_pc_10,
	F_pc_11,
	F_pc_12,
	F_pc_14,
	q_a_0,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_12,
	q_a_14,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	F_pc_2,
	q_a_8,
	q_a_10,
	q_a_17,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_5,
	F_pc_4,
	F_pc_3,
	q_a_9,
	q_a_6,
	F_pc_1,
	q_a_7,
	F_pc_0,
	readdata_0,
	q_b_0,
	readdata_22,
	d_writedata_22,
	readdata_23,
	d_writedata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_11,
	d_writedata_11,
	readdata_12,
	d_writedata_12,
	readdata_13,
	d_writedata_13,
	readdata_14,
	d_writedata_14,
	readdata_15,
	d_writedata_15,
	readdata_16,
	d_writedata_16,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_8,
	d_writedata_8,
	q_a_27,
	q_a_28,
	q_a_29,
	q_a_30,
	q_a_31,
	readdata_10,
	d_writedata_10,
	readdata_17,
	d_writedata_17,
	readdata_9,
	d_writedata_9,
	readdata_18,
	d_writedata_18,
	readdata_19,
	d_writedata_19,
	readdata_20,
	d_writedata_20,
	readdata_21,
	d_writedata_21,
	av_readdata_pre_16,
	readdata_6,
	readdata_7,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	readdata_27,
	readdata_28,
	readdata_29,
	readdata_30,
	readdata_31,
	av_readdata_pre_19,
	av_readdata_pre_18,
	av_readdata_pre_17,
	q_b_7,
	q_b_6,
	av_readdata_pre_20,
	av_readdata_pre_21,
	av_readdata_pre_22,
	Add1,
	Add11,
	Add12,
	Add13,
	Add14,
	Add15,
	Add16,
	nios2_gen2_0_data_master_waitrequest,
	d_writedata_0,
	r_sync_rst,
	mem_used_1,
	Equal2,
	Equal21,
	rst1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	d_write,
	write_accepted,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	always0,
	d_read,
	read_accepted,
	always2,
	av_waitrequest,
	always01,
	read_latency_shift_reg,
	saved_grant_0,
	waitrequest,
	mem_used_11,
	saved_grant_01,
	mem_used_12,
	Equal3,
	mem_used_13,
	av_waitrequest1,
	WideOr0,
	src0_valid,
	read_latency_shift_reg_0,
	WideOr1,
	av_waitrequest2,
	src1_valid,
	i_read,
	F_pc_13,
	src_valid,
	mem,
	src2_valid,
	src_valid1,
	hbreak_enabled,
	av_waitrequest3,
	src0_valid1,
	src_data_0,
	av_readdata_pre_221,
	src1_valid1,
	src1_valid2,
	src_data_22,
	av_readdata_pre_23,
	src_data_23,
	src_data_24,
	src_data_25,
	src_data_26,
	av_readdata_pre_11,
	av_readdata_pre_12,
	src_data_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	src_data_14,
	av_readdata_pre_15,
	av_readdata_pre_161,
	src_data_01,
	av_readdata_pre_1,
	src_data_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_8,
	src_data_8,
	av_readdata_pre_10,
	src_data_10,
	av_readdata_pre_171,
	src_data_17,
	av_readdata_pre_9,
	src_data_9,
	av_readdata_pre_181,
	av_readdata_pre_191,
	av_readdata_pre_201,
	av_readdata_pre_211,
	src_data_6,
	src_data_46,
	src_data_7,
	src_data_1,
	src_data_21,
	src_data_3,
	src_data_4,
	src_data_5,
	b_full,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_461,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	d_byteenable_0,
	src_data_32,
	ien_AF,
	read_0,
	readdata_01,
	av_readdata_pre_81,
	src_payload1,
	d_byteenable_2,
	src_data_34,
	src_payload2,
	d_writedata_24,
	src_payload3,
	d_byteenable_3,
	src_data_35,
	d_writedata_25,
	src_payload4,
	d_writedata_26,
	src_payload5,
	src_payload6,
	d_byteenable_1,
	src_data_33,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_data_27,
	src_data_28,
	src_data_29,
	src_data_30,
	src_data_31,
	src_payload18,
	src_payload19,
	av_readdata_pre_101,
	av_readdata_pre_91,
	src_payload20,
	src_payload21,
	src_payload22,
	av_readdata_pre_121,
	src_payload23,
	av_readdata_pre_131,
	src_payload24,
	av_readdata_pre_141,
	src_payload25,
	av_readdata_pre_151,
	src_payload26,
	d_writedata_6,
	src_payload27,
	d_writedata_7,
	src_payload28,
	ien_AE,
	readdata_110,
	readdata_210,
	readdata_32,
	readdata_41,
	readdata_51,
	b_non_empty,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	src_payload29,
	src_data_381,
	src_data_411,
	src_data_451,
	src_data_441,
	src_data_431,
	src_data_421,
	src_data_401,
	src_data_391,
	src_payload30,
	src_data_321,
	av_readdata_8,
	d_writedata_27,
	src_payload31,
	d_writedata_28,
	src_payload32,
	d_writedata_29,
	src_payload33,
	d_writedata_30,
	src_payload34,
	d_writedata_31,
	src_payload35,
	ac,
	av_readdata_9,
	b_full1,
	woverflow,
	rvalid,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_payload41,
	src_payload42,
	src_payload43,
	src_payload44,
	src_payload45,
	src_payload46,
	src_payload47,
	src_data_341,
	src_payload48,
	src_payload49,
	src_data_351,
	src_payload50,
	src_payload51,
	src_payload52,
	src_data_331,
	src_payload53,
	src_payload54,
	src_payload55,
	src_payload56,
	src_payload57,
	src_payload58,
	src_payload59,
	src_payload60,
	src_payload61,
	src_payload62,
	src_payload63,
	src_payload64,
	src_payload65,
	src_payload66,
	src_payload67,
	src_payload68,
	src_payload69,
	src_payload70,
	src_payload71,
	src_payload72,
	src_payload73,
	src_payload74,
	GND_port,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_7;
input 	W_alu_result_6;
input 	W_alu_result_5;
input 	W_alu_result_12;
input 	W_alu_result_13;
input 	W_alu_result_14;
input 	W_alu_result_15;
input 	W_alu_result_16;
input 	W_alu_result_3;
input 	W_alu_result_2;
input 	F_pc_9;
input 	F_pc_10;
input 	F_pc_11;
input 	F_pc_12;
input 	F_pc_14;
input 	q_a_0;
input 	q_a_22;
input 	q_a_23;
input 	q_a_24;
input 	q_a_25;
input 	q_a_26;
input 	q_a_12;
input 	q_a_14;
input 	q_a_1;
input 	q_a_2;
input 	q_a_3;
input 	q_a_4;
input 	q_a_5;
input 	F_pc_2;
input 	q_a_8;
input 	q_a_10;
input 	q_a_17;
input 	F_pc_8;
input 	F_pc_7;
input 	F_pc_6;
input 	F_pc_5;
input 	F_pc_4;
input 	F_pc_3;
input 	q_a_9;
input 	q_a_6;
input 	F_pc_1;
input 	q_a_7;
input 	F_pc_0;
input 	readdata_0;
input 	q_b_0;
input 	readdata_22;
input 	d_writedata_22;
input 	readdata_23;
input 	d_writedata_23;
input 	readdata_24;
input 	readdata_25;
input 	readdata_26;
input 	readdata_11;
input 	d_writedata_11;
input 	readdata_12;
input 	d_writedata_12;
input 	readdata_13;
input 	d_writedata_13;
input 	readdata_14;
input 	d_writedata_14;
input 	readdata_15;
input 	d_writedata_15;
input 	readdata_16;
input 	d_writedata_16;
input 	readdata_1;
input 	readdata_2;
input 	readdata_3;
input 	readdata_4;
input 	readdata_5;
input 	readdata_8;
input 	d_writedata_8;
input 	q_a_27;
input 	q_a_28;
input 	q_a_29;
input 	q_a_30;
input 	q_a_31;
input 	readdata_10;
input 	d_writedata_10;
input 	readdata_17;
input 	d_writedata_17;
input 	readdata_9;
input 	d_writedata_9;
input 	readdata_18;
input 	d_writedata_18;
input 	readdata_19;
input 	d_writedata_19;
input 	readdata_20;
input 	d_writedata_20;
input 	readdata_21;
input 	d_writedata_21;
output 	av_readdata_pre_16;
input 	readdata_6;
input 	readdata_7;
input 	q_b_1;
input 	q_b_2;
input 	q_b_3;
input 	q_b_4;
input 	q_b_5;
input 	readdata_27;
input 	readdata_28;
input 	readdata_29;
input 	readdata_30;
input 	readdata_31;
output 	av_readdata_pre_19;
output 	av_readdata_pre_18;
output 	av_readdata_pre_17;
input 	q_b_7;
input 	q_b_6;
output 	av_readdata_pre_20;
output 	av_readdata_pre_21;
output 	av_readdata_pre_22;
input 	Add1;
input 	Add11;
input 	Add12;
input 	Add13;
input 	Add14;
input 	Add15;
input 	Add16;
output 	nios2_gen2_0_data_master_waitrequest;
input 	d_writedata_0;
input 	r_sync_rst;
output 	mem_used_1;
output 	Equal2;
output 	Equal21;
input 	rst1;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	d_write;
output 	write_accepted;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	always0;
input 	d_read;
output 	read_accepted;
input 	always2;
output 	av_waitrequest;
input 	always01;
output 	read_latency_shift_reg;
output 	saved_grant_0;
input 	waitrequest;
output 	mem_used_11;
output 	saved_grant_01;
output 	mem_used_12;
output 	Equal3;
output 	mem_used_13;
input 	av_waitrequest1;
output 	WideOr0;
output 	src0_valid;
output 	read_latency_shift_reg_0;
output 	WideOr1;
input 	av_waitrequest2;
output 	src1_valid;
input 	i_read;
input 	F_pc_13;
output 	src_valid;
output 	mem;
output 	src2_valid;
output 	src_valid1;
input 	hbreak_enabled;
output 	av_waitrequest3;
output 	src0_valid1;
output 	src_data_0;
output 	av_readdata_pre_221;
output 	src1_valid1;
output 	src1_valid2;
output 	src_data_22;
output 	av_readdata_pre_23;
output 	src_data_23;
output 	src_data_24;
output 	src_data_25;
output 	src_data_26;
output 	av_readdata_pre_11;
output 	av_readdata_pre_12;
output 	src_data_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	src_data_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_161;
output 	src_data_01;
output 	av_readdata_pre_1;
output 	src_data_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_8;
output 	src_data_8;
output 	av_readdata_pre_10;
output 	src_data_10;
output 	av_readdata_pre_171;
output 	src_data_17;
output 	av_readdata_pre_9;
output 	src_data_9;
output 	av_readdata_pre_181;
output 	av_readdata_pre_191;
output 	av_readdata_pre_201;
output 	av_readdata_pre_211;
output 	src_data_6;
output 	src_data_46;
output 	src_data_7;
output 	src_data_1;
output 	src_data_21;
output 	src_data_3;
output 	src_data_4;
output 	src_data_5;
input 	b_full;
output 	src_payload;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_461;
output 	src_data_47;
output 	src_data_48;
output 	src_data_49;
output 	src_data_50;
input 	d_byteenable_0;
output 	src_data_32;
input 	ien_AF;
input 	read_0;
input 	readdata_01;
output 	av_readdata_pre_81;
output 	src_payload1;
input 	d_byteenable_2;
output 	src_data_34;
output 	src_payload2;
input 	d_writedata_24;
output 	src_payload3;
input 	d_byteenable_3;
output 	src_data_35;
input 	d_writedata_25;
output 	src_payload4;
input 	d_writedata_26;
output 	src_payload5;
output 	src_payload6;
input 	d_byteenable_1;
output 	src_data_33;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_data_27;
output 	src_data_28;
output 	src_data_29;
output 	src_data_30;
output 	src_data_31;
output 	src_payload18;
output 	src_payload19;
output 	av_readdata_pre_101;
output 	av_readdata_pre_91;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	av_readdata_pre_121;
output 	src_payload23;
output 	av_readdata_pre_131;
output 	src_payload24;
output 	av_readdata_pre_141;
output 	src_payload25;
output 	av_readdata_pre_151;
output 	src_payload26;
input 	d_writedata_6;
output 	src_payload27;
input 	d_writedata_7;
output 	src_payload28;
input 	ien_AE;
input 	readdata_110;
input 	readdata_210;
input 	readdata_32;
input 	readdata_41;
input 	readdata_51;
input 	b_non_empty;
input 	counter_reg_bit_1;
input 	counter_reg_bit_0;
input 	counter_reg_bit_5;
input 	counter_reg_bit_4;
input 	counter_reg_bit_3;
input 	counter_reg_bit_2;
output 	src_payload29;
output 	src_data_381;
output 	src_data_411;
output 	src_data_451;
output 	src_data_441;
output 	src_data_431;
output 	src_data_421;
output 	src_data_401;
output 	src_data_391;
output 	src_payload30;
output 	src_data_321;
input 	av_readdata_8;
input 	d_writedata_27;
output 	src_payload31;
input 	d_writedata_28;
output 	src_payload32;
input 	d_writedata_29;
output 	src_payload33;
input 	d_writedata_30;
output 	src_payload34;
input 	d_writedata_31;
output 	src_payload35;
input 	ac;
input 	av_readdata_9;
input 	b_full1;
input 	woverflow;
input 	rvalid;
output 	src_payload36;
output 	src_payload37;
output 	src_payload38;
output 	src_payload39;
output 	src_payload40;
output 	src_payload41;
output 	src_payload42;
output 	src_payload43;
output 	src_payload44;
output 	src_payload45;
output 	src_payload46;
output 	src_payload47;
output 	src_data_341;
output 	src_payload48;
output 	src_payload49;
output 	src_data_351;
output 	src_payload50;
output 	src_payload51;
output 	src_payload52;
output 	src_data_331;
output 	src_payload53;
output 	src_payload54;
output 	src_payload55;
output 	src_payload56;
output 	src_payload57;
output 	src_payload58;
output 	src_payload59;
output 	src_payload60;
output 	src_payload61;
output 	src_payload62;
output 	src_payload63;
output 	src_payload64;
output 	src_payload65;
output 	src_payload66;
output 	src_payload67;
output 	src_payload68;
output 	src_payload69;
output 	src_payload70;
output 	src_payload71;
output 	src_payload72;
output 	src_payload73;
output 	src_payload74;
input 	GND_port;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[0]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[1]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[2]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[3]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[4]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[5]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[7]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[6]~q ;
wire \pio_0_s1_translator|read_latency_shift_reg~0_combout ;
wire \pio_0_s1_agent|m0_write~0_combout ;
wire \pio_0_s1_translator|av_waitrequest_generated~0_combout ;
wire \pio_0_s1_translator|read_latency_shift_reg[0]~q ;
wire \pio_0_s1_agent|m0_write~1_combout ;
wire \router|Equal2~2_combout ;
wire \router|Equal1~0_combout ;
wire \cmd_demux|WideOr0~2_combout ;
wire \cmd_demux|sink_ready~0_combout ;
wire \onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem[0][56]~q ;
wire \nios2_gen2_0_debug_mem_slave_translator|read_latency_shift_reg[0]~q ;
wire \nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem[0][74]~q ;
wire \nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem[0][56]~q ;
wire \cmd_demux|WideOr0~4_combout ;
wire \cmd_demux|WideOr0~5_combout ;
wire \jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ;
wire \nios2_gen2_0_instruction_master_translator|read_accepted~q ;
wire \router_001|Equal1~0_combout ;
wire \cmd_demux_001|src0_valid~0_combout ;
wire \nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|write~0_combout ;
wire \cmd_mux_001|saved_grant[1]~q ;
wire \cmd_demux_001|src1_valid~0_combout ;
wire \onchip_memory2_0_s1_translator|read_latency_shift_reg~0_combout ;
wire \cmd_mux_002|saved_grant[1]~q ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem~0_combout ;
wire \cmd_demux|sink_ready~1_combout ;
wire \nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[0]~q ;
wire \pio_0_s1_translator|av_readdata_pre[0]~q ;
wire \nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[24]~q ;
wire \nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[25]~q ;
wire \nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[26]~q ;
wire \nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[2]~q ;
wire \nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[6]~q ;
wire \nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[7]~q ;
wire \pio_0_s1_translator|av_readdata_pre[1]~q ;
wire \pio_0_s1_translator|av_readdata_pre[2]~q ;
wire \pio_0_s1_translator|av_readdata_pre[3]~q ;
wire \pio_0_s1_translator|av_readdata_pre[4]~q ;
wire \pio_0_s1_translator|av_readdata_pre[5]~q ;
wire \nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[27]~q ;
wire \nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[28]~q ;
wire \nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[29]~q ;
wire \nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[30]~q ;
wire \nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[31]~q ;


niosLab2_niosLab2_mm_interconnect_0_rsp_mux_001 rsp_mux_001(
	.q_a_0(q_a_0),
	.q_a_22(q_a_22),
	.q_a_23(q_a_23),
	.q_a_24(q_a_24),
	.q_a_25(q_a_25),
	.q_a_26(q_a_26),
	.q_a_12(q_a_12),
	.q_a_14(q_a_14),
	.q_a_2(q_a_2),
	.q_a_8(q_a_8),
	.q_a_10(q_a_10),
	.q_a_17(q_a_17),
	.q_a_9(q_a_9),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.q_a_27(q_a_27),
	.q_a_28(q_a_28),
	.q_a_29(q_a_29),
	.q_a_30(q_a_30),
	.q_a_31(q_a_31),
	.av_readdata_pre_0(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_22(av_readdata_pre_221),
	.src1_valid(src1_valid1),
	.src1_valid1(src1_valid2),
	.src_data_22(src_data_22),
	.av_readdata_pre_23(av_readdata_pre_23),
	.src_data_23(src_data_23),
	.av_readdata_pre_24(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[24]~q ),
	.src_data_24(src_data_24),
	.av_readdata_pre_25(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[25]~q ),
	.src_data_25(src_data_25),
	.av_readdata_pre_26(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[26]~q ),
	.src_data_26(src_data_26),
	.av_readdata_pre_12(av_readdata_pre_12),
	.src_data_12(src_data_12),
	.av_readdata_pre_14(av_readdata_pre_14),
	.src_data_14(src_data_14),
	.src_data_0(src_data_01),
	.av_readdata_pre_2(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[2]~q ),
	.src_data_2(src_data_2),
	.av_readdata_pre_8(av_readdata_pre_8),
	.src_data_8(src_data_8),
	.av_readdata_pre_10(av_readdata_pre_10),
	.src_data_10(src_data_10),
	.av_readdata_pre_17(av_readdata_pre_171),
	.src_data_17(src_data_17),
	.av_readdata_pre_9(av_readdata_pre_9),
	.src_data_9(src_data_9),
	.av_readdata_pre_6(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[6]~q ),
	.src_data_6(src_data_6),
	.av_readdata_pre_7(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[7]~q ),
	.src_data_7(src_data_7),
	.av_readdata_pre_27(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[27]~q ),
	.src_data_27(src_data_27),
	.av_readdata_pre_28(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[28]~q ),
	.src_data_28(src_data_28),
	.av_readdata_pre_29(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[29]~q ),
	.src_data_29(src_data_29),
	.av_readdata_pre_30(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[30]~q ),
	.src_data_30(src_data_30),
	.av_readdata_pre_31(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[31]~q ),
	.src_data_31(src_data_31));

niosLab2_niosLab2_mm_interconnect_0_rsp_mux rsp_mux(
	.q_a_0(q_a_0),
	.av_readdata_pre_0(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.q_a_24(q_a_24),
	.q_a_25(q_a_25),
	.q_a_26(q_a_26),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.av_readdata_pre_1(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.q_a_27(q_a_27),
	.q_a_28(q_a_28),
	.q_a_29(q_a_29),
	.q_a_30(q_a_30),
	.q_a_31(q_a_31),
	.av_readdata_pre_7(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_6(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.read_latency_shift_reg_0(\pio_0_s1_translator|read_latency_shift_reg[0]~q ),
	.src0_valid(src0_valid),
	.read_latency_shift_reg_01(read_latency_shift_reg_0),
	.read_latency_shift_reg_02(\nios2_gen2_0_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem[0][56]~q ),
	.WideOr1(WideOr1),
	.src0_valid1(src0_valid1),
	.av_readdata_pre_01(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_02(\pio_0_s1_translator|av_readdata_pre[0]~q ),
	.src_data_0(src_data_0),
	.av_readdata_pre_24(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_25(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_26(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[26]~q ),
	.av_readdata_pre_11(av_readdata_pre_1),
	.av_readdata_pre_21(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_31(av_readdata_pre_3),
	.av_readdata_pre_41(av_readdata_pre_4),
	.av_readdata_pre_51(av_readdata_pre_5),
	.av_readdata_pre_61(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_71(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_12(\pio_0_s1_translator|av_readdata_pre[1]~q ),
	.src_data_1(src_data_1),
	.av_readdata_pre_22(\pio_0_s1_translator|av_readdata_pre[2]~q ),
	.src_data_2(src_data_21),
	.av_readdata_pre_32(\pio_0_s1_translator|av_readdata_pre[3]~q ),
	.src_data_3(src_data_3),
	.av_readdata_pre_42(\pio_0_s1_translator|av_readdata_pre[4]~q ),
	.src_data_4(src_data_4),
	.av_readdata_pre_52(\pio_0_s1_translator|av_readdata_pre[5]~q ),
	.src_data_5(src_data_5),
	.av_readdata_pre_27(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_28(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_29(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_30(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_311(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[31]~q ),
	.src_payload(src_payload20),
	.src_payload1(src_payload21),
	.src_payload2(src_payload36),
	.src_payload3(src_payload38),
	.src_payload4(src_payload39),
	.src_payload5(src_payload40),
	.src_payload6(src_payload41),
	.src_payload7(src_payload42),
	.src_payload8(src_payload43),
	.src_payload9(src_payload44));

niosLab2_niosLab2_mm_interconnect_0_cmd_demux_001_2 rsp_demux_002(
	.read_latency_shift_reg_0(\onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid(src0_valid),
	.src1_valid(src1_valid2));

niosLab2_niosLab2_mm_interconnect_0_cmd_demux_001_1 rsp_demux_001(
	.read_latency_shift_reg_0(\nios2_gen2_0_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid(src0_valid1),
	.src1_valid(src1_valid1));

niosLab2_niosLab2_mm_interconnect_0_cmd_mux_001_1 cmd_mux_002(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_3(W_alu_result_3),
	.W_alu_result_2(W_alu_result_2),
	.F_pc_9(F_pc_9),
	.F_pc_10(F_pc_10),
	.F_pc_11(F_pc_11),
	.F_pc_12(F_pc_12),
	.F_pc_2(F_pc_2),
	.F_pc_8(F_pc_8),
	.F_pc_7(F_pc_7),
	.F_pc_6(F_pc_6),
	.F_pc_5(F_pc_5),
	.F_pc_4(F_pc_4),
	.F_pc_3(F_pc_3),
	.F_pc_1(F_pc_1),
	.F_pc_0(F_pc_0),
	.d_writedata_22(d_writedata_22),
	.d_writedata_23(d_writedata_23),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.d_writedata_16(d_writedata_16),
	.d_writedata_8(d_writedata_8),
	.d_writedata_10(d_writedata_10),
	.d_writedata_17(d_writedata_17),
	.d_writedata_9(d_writedata_9),
	.d_writedata_18(d_writedata_18),
	.d_writedata_19(d_writedata_19),
	.d_writedata_20(d_writedata_20),
	.d_writedata_21(d_writedata_21),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.rst1(rst1),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.saved_grant_0(saved_grant_01),
	.i_read(i_read),
	.read_accepted(\nios2_gen2_0_instruction_master_translator|read_accepted~q ),
	.Equal1(\router_001|Equal1~0_combout ),
	.src2_valid(src2_valid),
	.src1_valid(\cmd_demux_001|src1_valid~0_combout ),
	.read_latency_shift_reg(\onchip_memory2_0_s1_translator|read_latency_shift_reg~0_combout ),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.src_valid(src_valid1),
	.src_payload(src_payload),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.src_data_40(src_data_40),
	.src_data_41(src_data_41),
	.src_data_42(src_data_42),
	.src_data_43(src_data_43),
	.src_data_44(src_data_44),
	.src_data_45(src_data_45),
	.src_data_46(src_data_461),
	.src_data_47(src_data_47),
	.src_data_48(src_data_48),
	.src_data_49(src_data_49),
	.src_data_50(src_data_50),
	.d_byteenable_0(d_byteenable_0),
	.src_data_32(src_data_32),
	.src_payload1(src_payload1),
	.d_byteenable_2(d_byteenable_2),
	.src_data_34(src_data_34),
	.src_payload2(src_payload2),
	.d_writedata_24(d_writedata_24),
	.src_payload3(src_payload3),
	.d_byteenable_3(d_byteenable_3),
	.src_data_35(src_data_35),
	.d_writedata_25(d_writedata_25),
	.src_payload4(src_payload4),
	.d_writedata_26(d_writedata_26),
	.src_payload5(src_payload5),
	.src_payload6(src_payload6),
	.d_byteenable_1(d_byteenable_1),
	.src_data_33(src_data_33),
	.src_payload7(src_payload7),
	.src_payload8(src_payload8),
	.src_payload9(src_payload9),
	.src_payload10(src_payload10),
	.src_payload11(src_payload11),
	.src_payload12(src_payload12),
	.src_payload13(src_payload13),
	.src_payload14(src_payload14),
	.src_payload15(src_payload15),
	.src_payload16(src_payload16),
	.src_payload17(src_payload17),
	.src_payload18(src_payload18),
	.src_payload19(src_payload19),
	.src_payload20(src_payload22),
	.src_payload21(src_payload23),
	.src_payload22(src_payload24),
	.src_payload23(src_payload25),
	.src_payload24(src_payload26),
	.d_writedata_6(d_writedata_6),
	.src_payload25(src_payload27),
	.d_writedata_7(d_writedata_7),
	.src_payload26(src_payload28),
	.d_writedata_27(d_writedata_27),
	.src_payload27(src_payload31),
	.d_writedata_28(d_writedata_28),
	.src_payload28(src_payload32),
	.d_writedata_29(d_writedata_29),
	.src_payload29(src_payload33),
	.d_writedata_30(d_writedata_30),
	.src_payload30(src_payload34),
	.d_writedata_31(d_writedata_31),
	.src_payload31(src_payload35),
	.clk_clk(clk_clk));

niosLab2_niosLab2_mm_interconnect_0_cmd_mux_001 cmd_mux_001(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_3(W_alu_result_3),
	.W_alu_result_2(W_alu_result_2),
	.F_pc_2(F_pc_2),
	.F_pc_8(F_pc_8),
	.F_pc_7(F_pc_7),
	.F_pc_6(F_pc_6),
	.F_pc_5(F_pc_5),
	.F_pc_4(F_pc_4),
	.F_pc_3(F_pc_3),
	.F_pc_1(F_pc_1),
	.F_pc_0(F_pc_0),
	.d_writedata_22(d_writedata_22),
	.d_writedata_23(d_writedata_23),
	.d_writedata_11(d_writedata_11),
	.d_writedata_12(d_writedata_12),
	.d_writedata_13(d_writedata_13),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.d_writedata_16(d_writedata_16),
	.d_writedata_8(d_writedata_8),
	.d_writedata_10(d_writedata_10),
	.d_writedata_17(d_writedata_17),
	.d_writedata_9(d_writedata_9),
	.d_writedata_18(d_writedata_18),
	.d_writedata_19(d_writedata_19),
	.d_writedata_20(d_writedata_20),
	.d_writedata_21(d_writedata_21),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.rst1(rst1),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.saved_grant_0(saved_grant_0),
	.src1_valid(src1_valid),
	.i_read(i_read),
	.read_accepted(\nios2_gen2_0_instruction_master_translator|read_accepted~q ),
	.Equal1(\router_001|Equal1~0_combout ),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ),
	.write(\nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.src_valid(src_valid),
	.hbreak_enabled(hbreak_enabled),
	.src_data_46(src_data_46),
	.d_byteenable_0(d_byteenable_0),
	.d_byteenable_2(d_byteenable_2),
	.d_writedata_24(d_writedata_24),
	.d_byteenable_3(d_byteenable_3),
	.d_writedata_25(d_writedata_25),
	.d_writedata_26(d_writedata_26),
	.d_byteenable_1(d_byteenable_1),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.src_payload(src_payload29),
	.src_data_38(src_data_381),
	.src_data_41(src_data_411),
	.src_data_45(src_data_451),
	.src_data_44(src_data_441),
	.src_data_43(src_data_431),
	.src_data_42(src_data_421),
	.src_data_40(src_data_401),
	.src_data_39(src_data_391),
	.src_payload1(src_payload30),
	.src_data_32(src_data_321),
	.d_writedata_27(d_writedata_27),
	.d_writedata_28(d_writedata_28),
	.d_writedata_29(d_writedata_29),
	.d_writedata_30(d_writedata_30),
	.d_writedata_31(d_writedata_31),
	.src_payload2(src_payload37),
	.src_payload3(src_payload45),
	.src_payload4(src_payload46),
	.src_payload5(src_payload47),
	.src_data_34(src_data_341),
	.src_payload6(src_payload48),
	.src_payload7(src_payload49),
	.src_data_35(src_data_351),
	.src_payload8(src_payload50),
	.src_payload9(src_payload51),
	.src_payload10(src_payload52),
	.src_data_33(src_data_331),
	.src_payload11(src_payload53),
	.src_payload12(src_payload54),
	.src_payload13(src_payload55),
	.src_payload14(src_payload56),
	.src_payload15(src_payload57),
	.src_payload16(src_payload58),
	.src_payload17(src_payload59),
	.src_payload18(src_payload60),
	.src_payload19(src_payload61),
	.src_payload20(src_payload62),
	.src_payload21(src_payload63),
	.src_payload22(src_payload64),
	.src_payload23(src_payload65),
	.src_payload24(src_payload66),
	.src_payload25(src_payload67),
	.src_payload26(src_payload68),
	.src_payload27(src_payload69),
	.src_payload28(src_payload70),
	.src_payload29(src_payload71),
	.src_payload30(src_payload72),
	.src_payload31(src_payload73),
	.src_payload32(src_payload74),
	.clk_clk(clk_clk));

niosLab2_niosLab2_mm_interconnect_0_cmd_demux_001 cmd_demux_001(
	.rst1(rst1),
	.i_read(i_read),
	.read_accepted(\nios2_gen2_0_instruction_master_translator|read_accepted~q ),
	.Equal1(\router_001|Equal1~0_combout ),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ),
	.src1_valid(\cmd_demux_001|src1_valid~0_combout ));

niosLab2_niosLab2_mm_interconnect_0_cmd_demux cmd_demux(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_3(W_alu_result_3),
	.Equal2(Equal2),
	.Equal21(Equal21),
	.rst1(rst1),
	.av_waitrequest_generated(\pio_0_s1_translator|av_waitrequest_generated~0_combout ),
	.always0(always01),
	.Equal1(\router|Equal1~0_combout ),
	.saved_grant_0(saved_grant_0),
	.waitrequest(waitrequest),
	.mem_used_1(mem_used_11),
	.saved_grant_01(saved_grant_01),
	.mem_used_11(mem_used_12),
	.WideOr0(\cmd_demux|WideOr0~2_combout ),
	.Equal3(Equal3),
	.mem_used_12(mem_used_13),
	.av_waitrequest(av_waitrequest1),
	.sink_ready(\cmd_demux|sink_ready~0_combout ),
	.WideOr01(WideOr0),
	.WideOr02(\cmd_demux|WideOr0~4_combout ),
	.WideOr03(\cmd_demux|WideOr0~5_combout ),
	.av_waitrequest1(av_waitrequest2),
	.src1_valid(src1_valid),
	.src2_valid(src2_valid),
	.sink_ready1(\cmd_demux|sink_ready~1_combout ));

niosLab2_niosLab2_mm_interconnect_0_router_001 router_001(
	.F_pc_9(F_pc_9),
	.F_pc_10(F_pc_10),
	.F_pc_11(F_pc_11),
	.F_pc_12(F_pc_12),
	.F_pc_14(F_pc_14),
	.F_pc_13(F_pc_13),
	.Equal1(\router_001|Equal1~0_combout ));

niosLab2_niosLab2_mm_interconnect_0_router router(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_16(W_alu_result_16),
	.W_alu_result_3(W_alu_result_3),
	.Equal2(Equal2),
	.Equal21(Equal21),
	.Equal22(\router|Equal2~2_combout ),
	.Equal1(\router|Equal1~0_combout ),
	.Equal3(Equal3));

niosLab2_altera_merlin_master_translator_1 nios2_gen2_0_instruction_master_translator(
	.reset(r_sync_rst),
	.rst1(rst1),
	.mem_used_1(mem_used_12),
	.i_read(i_read),
	.read_accepted1(\nios2_gen2_0_instruction_master_translator|read_accepted~q ),
	.Equal1(\router_001|Equal1~0_combout ),
	.write(\nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.saved_grant_11(\cmd_mux_002|saved_grant[1]~q ),
	.src1_valid(src1_valid1),
	.src1_valid1(src1_valid2),
	.clk(clk_clk));

niosLab2_altera_merlin_master_translator nios2_gen2_0_data_master_translator(
	.av_waitrequest(nios2_gen2_0_data_master_waitrequest),
	.reset(r_sync_rst),
	.rst1(rst1),
	.d_write(d_write),
	.write_accepted1(write_accepted),
	.d_read(d_read),
	.read_accepted1(read_accepted),
	.read_latency_shift_reg(\pio_0_s1_translator|read_latency_shift_reg~0_combout ),
	.always2(always2),
	.av_waitrequest_generated(\pio_0_s1_translator|av_waitrequest_generated~0_combout ),
	.av_waitrequest1(av_waitrequest),
	.always0(always01),
	.read_latency_shift_reg1(read_latency_shift_reg),
	.WideOr0(\cmd_demux|WideOr0~2_combout ),
	.sink_ready(\cmd_demux|sink_ready~0_combout ),
	.WideOr01(WideOr0),
	.src0_valid(src0_valid),
	.WideOr1(WideOr1),
	.WideOr02(\cmd_demux|WideOr0~4_combout ),
	.WideOr03(\cmd_demux|WideOr0~5_combout ),
	.read_latency_shift_reg2(\jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ),
	.av_waitrequest2(av_waitrequest3),
	.clk(clk_clk));

niosLab2_altera_merlin_slave_translator_2 onchip_memory2_0_s1_translator(
	.reset(r_sync_rst),
	.rst1(rst1),
	.saved_grant_0(saved_grant_01),
	.mem_used_1(mem_used_12),
	.read_latency_shift_reg_0(\onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ),
	.src2_valid(src2_valid),
	.read_latency_shift_reg(\onchip_memory2_0_s1_translator|read_latency_shift_reg~0_combout ),
	.src_valid(src_valid1),
	.mem(\onchip_memory2_0_s1_agent_rsp_fifo|mem~0_combout ),
	.clk(clk_clk));

niosLab2_altera_merlin_slave_translator_1 nios2_gen2_0_debug_mem_slave_translator(
	.av_readdata({readdata_31,readdata_30,readdata_29,readdata_28,readdata_27,readdata_26,readdata_25,readdata_24,readdata_23,readdata_22,readdata_21,readdata_20,readdata_19,readdata_18,readdata_17,readdata_16,readdata_15,readdata_14,readdata_13,readdata_12,readdata_11,readdata_10,readdata_9,
readdata_8,readdata_7,readdata_6,readdata_5,readdata_4,readdata_3,readdata_2,readdata_1,readdata_0}),
	.reset(r_sync_rst),
	.rst1(rst1),
	.saved_grant_0(saved_grant_0),
	.read_latency_shift_reg_0(\nios2_gen2_0_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.src1_valid(src1_valid),
	.write(\nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.src_valid(src_valid),
	.mem(mem),
	.av_readdata_pre_0(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_22(av_readdata_pre_221),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_24(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_25(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_26(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[26]~q ),
	.av_readdata_pre_11(av_readdata_pre_11),
	.av_readdata_pre_12(av_readdata_pre_12),
	.av_readdata_pre_13(av_readdata_pre_13),
	.av_readdata_pre_14(av_readdata_pre_14),
	.av_readdata_pre_15(av_readdata_pre_15),
	.av_readdata_pre_16(av_readdata_pre_161),
	.av_readdata_pre_1(av_readdata_pre_1),
	.av_readdata_pre_2(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(av_readdata_pre_3),
	.av_readdata_pre_4(av_readdata_pre_4),
	.av_readdata_pre_5(av_readdata_pre_5),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_17(av_readdata_pre_171),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_18(av_readdata_pre_181),
	.av_readdata_pre_19(av_readdata_pre_191),
	.av_readdata_pre_20(av_readdata_pre_201),
	.av_readdata_pre_21(av_readdata_pre_211),
	.av_readdata_pre_6(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_27(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_28(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_29(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_30(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_31(\nios2_gen2_0_debug_mem_slave_translator|av_readdata_pre[31]~q ),
	.clk(clk_clk));

niosLab2_altera_merlin_slave_translator jtag_uart_0_avalon_jtag_slave_translator(
	.av_readdata_pre_0(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.q_b_0(q_b_0),
	.av_readdata_pre_7(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_6(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_16(av_readdata_pre_16),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.av_readdata_pre_19(av_readdata_pre_19),
	.av_readdata_pre_18(av_readdata_pre_18),
	.av_readdata_pre_17(av_readdata_pre_17),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.av_readdata_pre_20(av_readdata_pre_20),
	.av_readdata_pre_21(av_readdata_pre_21),
	.av_readdata_pre_22(av_readdata_pre_22),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Add16,Add15,Add14,Add11,Add12,Add13,Add1,rvalid,woverflow,gnd,b_non_empty,gnd,ac,av_readdata_9,av_readdata_8,GND_port,GND_port,GND_port,GND_port,GND_port,GND_port,ien_AE,ien_AF}),
	.reset(r_sync_rst),
	.rst1(rst1),
	.d_read(d_read),
	.read_accepted(read_accepted),
	.sink_ready(\cmd_demux|sink_ready~0_combout ),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.read_latency_shift_reg(\jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ),
	.b_full(b_full),
	.read_0(read_0),
	.av_readdata_pre_8(av_readdata_pre_81),
	.av_readdata_pre_10(av_readdata_pre_101),
	.av_readdata_pre_9(av_readdata_pre_91),
	.av_readdata_pre_12(av_readdata_pre_121),
	.av_readdata_pre_13(av_readdata_pre_131),
	.av_readdata_pre_14(av_readdata_pre_141),
	.av_readdata_pre_15(av_readdata_pre_151),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.b_full1(b_full1),
	.clk(clk_clk));

niosLab2_altera_avalon_sc_fifo_3 pio_0_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.mem_used_1(mem_used_1),
	.always0(always0),
	.read_latency_shift_reg(\pio_0_s1_translator|read_latency_shift_reg~0_combout ),
	.av_waitrequest_generated(\pio_0_s1_translator|av_waitrequest_generated~0_combout ),
	.read_latency_shift_reg_0(\pio_0_s1_translator|read_latency_shift_reg[0]~q ),
	.always01(always01),
	.clk(clk_clk));

niosLab2_altera_merlin_slave_agent_3 pio_0_s1_agent(
	.W_alu_result_4(W_alu_result_4),
	.mem_used_1(mem_used_1),
	.Equal2(Equal2),
	.Equal21(Equal21),
	.rst1(rst1),
	.d_write(d_write),
	.write_accepted(write_accepted),
	.d_read(d_read),
	.read_accepted(read_accepted),
	.m0_write(\pio_0_s1_agent|m0_write~0_combout ),
	.m0_write1(\pio_0_s1_agent|m0_write~1_combout ));

niosLab2_altera_avalon_sc_fifo_2 onchip_memory2_0_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.rst1(rst1),
	.read_latency_shift_reg(\pio_0_s1_translator|read_latency_shift_reg~0_combout ),
	.saved_grant_0(saved_grant_01),
	.mem_used_1(mem_used_12),
	.read_latency_shift_reg_0(\onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][56]~q ),
	.i_read(i_read),
	.read_accepted(\nios2_gen2_0_instruction_master_translator|read_accepted~q ),
	.src2_valid(src2_valid),
	.read_latency_shift_reg1(\onchip_memory2_0_s1_translator|read_latency_shift_reg~0_combout ),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.src_valid(src_valid1),
	.mem(\onchip_memory2_0_s1_agent_rsp_fifo|mem~0_combout ),
	.clk(clk_clk));

niosLab2_altera_avalon_sc_fifo_1 nios2_gen2_0_debug_mem_slave_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg(\pio_0_s1_translator|read_latency_shift_reg~0_combout ),
	.saved_grant_0(saved_grant_0),
	.waitrequest(waitrequest),
	.mem_used_1(mem_used_11),
	.read_latency_shift_reg_0(\nios2_gen2_0_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|mem[0][56]~q ),
	.src1_valid(src1_valid),
	.i_read(i_read),
	.read_accepted(\nios2_gen2_0_instruction_master_translator|read_accepted~q ),
	.write(\nios2_gen2_0_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.src_valid(src_valid),
	.mem(mem),
	.clk(clk_clk));

niosLab2_altera_avalon_sc_fifo jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo(
	.reset(r_sync_rst),
	.mem_used_1(mem_used_13),
	.sink_ready(\cmd_demux|sink_ready~0_combout ),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.read_latency_shift_reg(\jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ),
	.sink_ready1(\cmd_demux|sink_ready~1_combout ),
	.clk(clk_clk));

niosLab2_altera_merlin_slave_translator_3 pio_0_s1_translator(
	.W_alu_result_4(W_alu_result_4),
	.reset(r_sync_rst),
	.Equal2(Equal2),
	.Equal21(Equal21),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.d_read(d_read),
	.read_accepted(read_accepted),
	.read_latency_shift_reg(\pio_0_s1_translator|read_latency_shift_reg~0_combout ),
	.always2(always2),
	.m0_write(\pio_0_s1_agent|m0_write~0_combout ),
	.av_waitrequest_generated(\pio_0_s1_translator|av_waitrequest_generated~0_combout ),
	.read_latency_shift_reg_0(\pio_0_s1_translator|read_latency_shift_reg[0]~q ),
	.m0_write1(\pio_0_s1_agent|m0_write~1_combout ),
	.Equal22(\router|Equal2~2_combout ),
	.always0(always01),
	.read_latency_shift_reg1(read_latency_shift_reg),
	.av_readdata_pre_0(\pio_0_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\pio_0_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\pio_0_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\pio_0_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\pio_0_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\pio_0_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_51,readdata_41,readdata_32,readdata_210,readdata_110,readdata_01}),
	.clk(clk_clk));

endmodule

module niosLab2_altera_avalon_sc_fifo (
	reset,
	mem_used_1,
	sink_ready,
	read_latency_shift_reg_0,
	read_latency_shift_reg,
	sink_ready1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	mem_used_1;
input 	sink_ready;
input 	read_latency_shift_reg_0;
input 	read_latency_shift_reg;
input 	sink_ready1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!sink_ready),
	.datac(!read_latency_shift_reg_0),
	.datad(!read_latency_shift_reg),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!sink_ready1),
	.datac(!read_latency_shift_reg_0),
	.datad(!read_latency_shift_reg),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hF3FF77FFF3FF77FF;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module niosLab2_altera_avalon_sc_fifo_1 (
	reset,
	read_latency_shift_reg,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src1_valid,
	i_read,
	read_accepted,
	write,
	saved_grant_1,
	src_valid,
	mem,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg;
input 	saved_grant_0;
input 	waitrequest;
output 	mem_used_1;
input 	read_latency_shift_reg_0;
output 	mem_74_0;
output 	mem_56_0;
input 	src1_valid;
input 	i_read;
input 	read_accepted;
output 	write;
input 	saved_grant_1;
input 	src_valid;
output 	mem;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~4_combout ;
wire \mem_used[0]~5_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;
wire \mem_used[1]~3_combout ;
wire \mem[1][74]~q ;
wire \mem~1_combout ;
wire \mem[1][56]~q ;
wire \mem~2_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][56] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_56_0),
	.prn(vcc));
defparam \mem[0][56] .is_wysiwyg = "true";
defparam \mem[0][56] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!waitrequest),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem~0 (
	.dataa(!read_latency_shift_reg),
	.datab(!saved_grant_0),
	.datac(!i_read),
	.datad(!read_accepted),
	.datae(!saved_grant_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(mem),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~4 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~4 .extended_lut = "off";
defparam \mem_used[0]~4 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \mem_used[0]~4 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~5 (
	.dataa(!saved_grant_0),
	.datab(!write),
	.datac(!src1_valid),
	.datad(!src_valid),
	.datae(!mem),
	.dataf(!\mem_used[0]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~5 .extended_lut = "off";
defparam \mem_used[0]~5 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \mem_used[0]~5 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \mem_used[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \mem_used[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~2 (
	.dataa(!waitrequest),
	.datab(!\mem_used[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~2 .extended_lut = "off";
defparam \mem_used[1]~2 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \mem_used[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~3 (
	.dataa(!saved_grant_0),
	.datab(!src1_valid),
	.datac(!src_valid),
	.datad(!mem),
	.datae(!\mem_used[1]~0_combout ),
	.dataf(!\mem_used[1]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~3 .extended_lut = "off";
defparam \mem_used[1]~3 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \mem_used[1]~3 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!saved_grant_1),
	.datac(!\mem[1][74]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][56] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][56]~q ),
	.prn(vcc));
defparam \mem[1][56] .is_wysiwyg = "true";
defparam \mem[1][56] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!mem),
	.datac(!\mem[1][56]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

endmodule

module niosLab2_altera_avalon_sc_fifo_2 (
	reset,
	rst1,
	read_latency_shift_reg,
	saved_grant_0,
	mem_used_1,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	i_read,
	read_accepted,
	src2_valid,
	read_latency_shift_reg1,
	saved_grant_1,
	src_valid,
	mem,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	rst1;
input 	read_latency_shift_reg;
input 	saved_grant_0;
output 	mem_used_1;
input 	read_latency_shift_reg_0;
output 	mem_74_0;
output 	mem_56_0;
input 	i_read;
input 	read_accepted;
input 	src2_valid;
input 	read_latency_shift_reg1;
input 	saved_grant_1;
input 	src_valid;
output 	mem;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~4_combout ;
wire \mem_used[0]~5_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;
wire \mem_used[1]~3_combout ;
wire \mem[1][74]~q ;
wire \mem~1_combout ;
wire \mem[1][56]~q ;
wire \mem~2_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][56] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_56_0),
	.prn(vcc));
defparam \mem[0][56] .is_wysiwyg = "true";
defparam \mem[0][56] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!read_latency_shift_reg),
	.datab(!saved_grant_0),
	.datac(!i_read),
	.datad(!read_accepted),
	.datae(!saved_grant_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(mem),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~4 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~4 .extended_lut = "off";
defparam \mem_used[0]~4 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \mem_used[0]~4 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~5 (
	.dataa(!saved_grant_0),
	.datab(!read_latency_shift_reg1),
	.datac(!src2_valid),
	.datad(!src_valid),
	.datae(!mem),
	.dataf(!\mem_used[0]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~5 .extended_lut = "off";
defparam \mem_used[0]~5 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \mem_used[0]~5 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \mem_used[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \mem_used[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~2 (
	.dataa(!rst1),
	.datab(!\mem_used[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~2 .extended_lut = "off";
defparam \mem_used[1]~2 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \mem_used[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~3 (
	.dataa(!saved_grant_0),
	.datab(!src2_valid),
	.datac(!src_valid),
	.datad(!mem),
	.datae(!\mem_used[1]~0_combout ),
	.dataf(!\mem_used[1]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~3 .extended_lut = "off";
defparam \mem_used[1]~3 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \mem_used[1]~3 .shared_arith = "off";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!saved_grant_1),
	.datac(!\mem[1][74]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][56] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][56]~q ),
	.prn(vcc));
defparam \mem[1][56] .is_wysiwyg = "true";
defparam \mem[1][56] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!mem),
	.datac(!\mem[1][56]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

endmodule

module niosLab2_altera_avalon_sc_fifo_3 (
	reset,
	mem_used_1,
	always0,
	read_latency_shift_reg,
	av_waitrequest_generated,
	read_latency_shift_reg_0,
	always01,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	mem_used_1;
input 	always0;
input 	read_latency_shift_reg;
input 	av_waitrequest_generated;
input 	read_latency_shift_reg_0;
input 	always01;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!always01),
	.datac(!read_latency_shift_reg),
	.datad(!av_waitrequest_generated),
	.datae(!read_latency_shift_reg_0),
	.dataf(!\mem_used[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!always0),
	.datac(!read_latency_shift_reg),
	.datad(!av_waitrequest_generated),
	.datae(!read_latency_shift_reg_0),
	.dataf(!\mem_used[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hFFFF3FFF7FFF7FFF;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module niosLab2_altera_merlin_master_translator (
	av_waitrequest,
	reset,
	rst1,
	d_write,
	write_accepted1,
	d_read,
	read_accepted1,
	read_latency_shift_reg,
	always2,
	av_waitrequest_generated,
	av_waitrequest1,
	always0,
	read_latency_shift_reg1,
	WideOr0,
	sink_ready,
	WideOr01,
	src0_valid,
	WideOr1,
	WideOr02,
	WideOr03,
	read_latency_shift_reg2,
	av_waitrequest2,
	clk)/* synthesis synthesis_greybox=1 */;
output 	av_waitrequest;
input 	reset;
input 	rst1;
input 	d_write;
output 	write_accepted1;
input 	d_read;
output 	read_accepted1;
input 	read_latency_shift_reg;
input 	always2;
input 	av_waitrequest_generated;
output 	av_waitrequest1;
input 	always0;
input 	read_latency_shift_reg1;
input 	WideOr0;
input 	sink_ready;
input 	WideOr01;
input 	src0_valid;
input 	WideOr1;
input 	WideOr02;
input 	WideOr03;
input 	read_latency_shift_reg2;
output 	av_waitrequest2;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \end_begintransfer~0_combout ;
wire \end_begintransfer~q ;
wire \write_accepted~0_combout ;
wire \read_accepted~0_combout ;
wire \read_accepted~1_combout ;


cyclonev_lcell_comb \av_waitrequest~2 (
	.dataa(!write_accepted1),
	.datab(!d_write),
	.datac(!WideOr1),
	.datad(!rst1),
	.datae(!d_read),
	.dataf(!src0_valid),
	.datag(!\end_begintransfer~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest~2 .extended_lut = "on";
defparam \av_waitrequest~2 .lut_mask = 64'h7FFFF7FF7FFFF7FF;
defparam \av_waitrequest~2 .shared_arith = "off";

dffeas write_accepted(
	.clk(clk),
	.d(\write_accepted~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(write_accepted1),
	.prn(vcc));
defparam write_accepted.is_wysiwyg = "true";
defparam write_accepted.power_up = "low";

dffeas read_accepted(
	.clk(clk),
	.d(\read_accepted~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_accepted1),
	.prn(vcc));
defparam read_accepted.is_wysiwyg = "true";
defparam read_accepted.power_up = "low";

cyclonev_lcell_comb \av_waitrequest~0 (
	.dataa(!write_accepted1),
	.datab(!d_read),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest1),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest~0 .extended_lut = "off";
defparam \av_waitrequest~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \av_waitrequest~0 .shared_arith = "off";

cyclonev_lcell_comb \av_waitrequest~1 (
	.dataa(!always0),
	.datab(!av_waitrequest_generated),
	.datac(!av_waitrequest1),
	.datad(!WideOr02),
	.datae(!WideOr0),
	.dataf(!sink_ready),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest2),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest~1 .extended_lut = "off";
defparam \av_waitrequest~1 .lut_mask = 64'hFFFFFFFFFFEFFFFF;
defparam \av_waitrequest~1 .shared_arith = "off";

cyclonev_lcell_comb \end_begintransfer~0 (
	.dataa(!rst1),
	.datab(!always2),
	.datac(!read_latency_shift_reg),
	.datad(!\end_begintransfer~q ),
	.datae(!read_latency_shift_reg1),
	.dataf(!WideOr01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\end_begintransfer~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \end_begintransfer~0 .extended_lut = "off";
defparam \end_begintransfer~0 .lut_mask = 64'hFFFFBFFFFFFFFFFF;
defparam \end_begintransfer~0 .shared_arith = "off";

dffeas end_begintransfer(
	.clk(clk),
	.d(\end_begintransfer~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\end_begintransfer~q ),
	.prn(vcc));
defparam end_begintransfer.is_wysiwyg = "true";
defparam end_begintransfer.power_up = "low";

cyclonev_lcell_comb \write_accepted~0 (
	.dataa(!rst1),
	.datab(!d_write),
	.datac(!write_accepted1),
	.datad(gnd),
	.datae(!WideOr03),
	.dataf(!av_waitrequest),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_accepted~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_accepted~0 .extended_lut = "off";
defparam \write_accepted~0 .lut_mask = 64'hFFFF7F7FFFFFFFFF;
defparam \write_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \read_accepted~0 (
	.dataa(!read_accepted1),
	.datab(!src0_valid),
	.datac(!WideOr1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_accepted~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_accepted~0 .extended_lut = "off";
defparam \read_accepted~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \read_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \read_accepted~1 (
	.dataa(gnd),
	.datab(!read_latency_shift_reg1),
	.datac(!WideOr01),
	.datad(!av_waitrequest),
	.datae(!\read_accepted~0_combout ),
	.dataf(!read_latency_shift_reg2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_accepted~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_accepted~1 .extended_lut = "off";
defparam \read_accepted~1 .lut_mask = 64'hF3FFFFFFFFFFFFFF;
defparam \read_accepted~1 .shared_arith = "off";

endmodule

module niosLab2_altera_merlin_master_translator_1 (
	reset,
	rst1,
	mem_used_1,
	i_read,
	read_accepted1,
	Equal1,
	write,
	saved_grant_1,
	saved_grant_11,
	src1_valid,
	src1_valid1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	rst1;
input 	mem_used_1;
input 	i_read;
output 	read_accepted1;
input 	Equal1;
input 	write;
input 	saved_grant_1;
input 	saved_grant_11;
input 	src1_valid;
input 	src1_valid1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_accepted~0_combout ;
wire \read_accepted~1_combout ;


dffeas read_accepted(
	.clk(clk),
	.d(\read_accepted~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_accepted1),
	.prn(vcc));
defparam read_accepted.is_wysiwyg = "true";
defparam read_accepted.power_up = "low";

cyclonev_lcell_comb \read_accepted~0 (
	.dataa(!write),
	.datab(!mem_used_1),
	.datac(!Equal1),
	.datad(!saved_grant_1),
	.datae(!saved_grant_11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_accepted~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_accepted~0 .extended_lut = "off";
defparam \read_accepted~0 .lut_mask = 64'hC5FFFFFFC5FFFFFF;
defparam \read_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \read_accepted~1 (
	.dataa(!rst1),
	.datab(!i_read),
	.datac(!read_accepted1),
	.datad(!src1_valid),
	.datae(!src1_valid1),
	.dataf(!\read_accepted~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_accepted~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_accepted~1 .extended_lut = "off";
defparam \read_accepted~1 .lut_mask = 64'hFFFFFFDFFFFFFFFF;
defparam \read_accepted~1 .shared_arith = "off";

endmodule

module niosLab2_altera_merlin_slave_agent_3 (
	W_alu_result_4,
	mem_used_1,
	Equal2,
	Equal21,
	rst1,
	d_write,
	write_accepted,
	d_read,
	read_accepted,
	m0_write,
	m0_write1)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	mem_used_1;
input 	Equal2;
input 	Equal21;
input 	rst1;
input 	d_write;
input 	write_accepted;
input 	d_read;
input 	read_accepted;
output 	m0_write;
output 	m0_write1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!mem_used_1),
	.datab(!rst1),
	.datac(!d_write),
	.datad(!write_accepted),
	.datae(!d_read),
	.dataf(!read_accepted),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hFFFFFFFFFFBFFFFF;
defparam \m0_write~0 .shared_arith = "off";

cyclonev_lcell_comb \m0_write~1 (
	.dataa(!W_alu_result_4),
	.datab(!Equal2),
	.datac(!Equal21),
	.datad(!m0_write),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~1 .extended_lut = "off";
defparam \m0_write~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \m0_write~1 .shared_arith = "off";

endmodule

module niosLab2_altera_merlin_slave_translator (
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	q_b_0,
	av_readdata_pre_7,
	av_readdata_pre_6,
	av_readdata_pre_16,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	av_readdata_pre_19,
	av_readdata_pre_18,
	av_readdata_pre_17,
	q_b_7,
	q_b_6,
	av_readdata_pre_20,
	av_readdata_pre_21,
	av_readdata_pre_22,
	av_readdata,
	reset,
	rst1,
	d_read,
	read_accepted,
	sink_ready,
	read_latency_shift_reg_0,
	read_latency_shift_reg,
	b_full,
	read_0,
	av_readdata_pre_8,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	b_full1,
	clk)/* synthesis synthesis_greybox=1 */;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
input 	q_b_0;
output 	av_readdata_pre_7;
output 	av_readdata_pre_6;
output 	av_readdata_pre_16;
input 	q_b_1;
input 	q_b_2;
input 	q_b_3;
input 	q_b_4;
input 	q_b_5;
output 	av_readdata_pre_19;
output 	av_readdata_pre_18;
output 	av_readdata_pre_17;
input 	q_b_7;
input 	q_b_6;
output 	av_readdata_pre_20;
output 	av_readdata_pre_21;
output 	av_readdata_pre_22;
input 	[31:0] av_readdata;
input 	reset;
input 	rst1;
input 	d_read;
input 	read_accepted;
input 	sink_ready;
output 	read_latency_shift_reg_0;
output 	read_latency_shift_reg;
input 	b_full;
input 	read_0;
output 	av_readdata_pre_8;
output 	av_readdata_pre_10;
output 	av_readdata_pre_9;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
input 	counter_reg_bit_1;
input 	counter_reg_bit_0;
input 	counter_reg_bit_5;
input 	counter_reg_bit_4;
input 	counter_reg_bit_3;
input 	counter_reg_bit_2;
input 	b_full1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~1_combout ;
wire \av_readdata_pre[13]~0_combout ;


dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(q_b_0),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(q_b_1),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(q_b_2),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(q_b_3),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(q_b_4),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(q_b_5),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(q_b_7),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(q_b_6),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(counter_reg_bit_0),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(counter_reg_bit_3),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(counter_reg_bit_2),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(counter_reg_bit_1),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(counter_reg_bit_4),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(counter_reg_bit_5),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(b_full),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!rst1),
	.datab(!d_read),
	.datac(!read_accepted),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(\av_readdata_pre[13]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!sink_ready),
	.datab(!read_latency_shift_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h7777777777777777;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \av_readdata_pre[13]~0 (
	.dataa(!b_full1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_readdata_pre[13]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdata_pre[13]~0 .extended_lut = "off";
defparam \av_readdata_pre[13]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \av_readdata_pre[13]~0 .shared_arith = "off";

endmodule

module niosLab2_altera_merlin_slave_translator_1 (
	av_readdata,
	reset,
	rst1,
	saved_grant_0,
	read_latency_shift_reg_0,
	src1_valid,
	write,
	src_valid,
	mem,
	av_readdata_pre_0,
	av_readdata_pre_22,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_16,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_8,
	av_readdata_pre_10,
	av_readdata_pre_17,
	av_readdata_pre_9,
	av_readdata_pre_18,
	av_readdata_pre_19,
	av_readdata_pre_20,
	av_readdata_pre_21,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_27,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_30,
	av_readdata_pre_31,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	reset;
input 	rst1;
input 	saved_grant_0;
output 	read_latency_shift_reg_0;
input 	src1_valid;
input 	write;
input 	src_valid;
input 	mem;
output 	av_readdata_pre_0;
output 	av_readdata_pre_22;
output 	av_readdata_pre_23;
output 	av_readdata_pre_24;
output 	av_readdata_pre_25;
output 	av_readdata_pre_26;
output 	av_readdata_pre_11;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_16;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_8;
output 	av_readdata_pre_10;
output 	av_readdata_pre_17;
output 	av_readdata_pre_9;
output 	av_readdata_pre_18;
output 	av_readdata_pre_19;
output 	av_readdata_pre_20;
output 	av_readdata_pre_21;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_27;
output 	av_readdata_pre_28;
output 	av_readdata_pre_29;
output 	av_readdata_pre_30;
output 	av_readdata_pre_31;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!rst1),
	.datab(!saved_grant_0),
	.datac(!write),
	.datad(!src1_valid),
	.datae(!src_valid),
	.dataf(!mem),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

endmodule

module niosLab2_altera_merlin_slave_translator_2 (
	reset,
	rst1,
	saved_grant_0,
	mem_used_1,
	read_latency_shift_reg_0,
	src2_valid,
	read_latency_shift_reg,
	src_valid,
	mem,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	rst1;
input 	saved_grant_0;
input 	mem_used_1;
output 	read_latency_shift_reg_0;
input 	src2_valid;
output 	read_latency_shift_reg;
input 	src_valid;
input 	mem;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~1_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!rst1),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!saved_grant_0),
	.datab(!read_latency_shift_reg),
	.datac(!src2_valid),
	.datad(!src_valid),
	.datae(!mem),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module niosLab2_altera_merlin_slave_translator_3 (
	W_alu_result_4,
	reset,
	Equal2,
	Equal21,
	wait_latency_counter_1,
	wait_latency_counter_0,
	d_read,
	read_accepted,
	read_latency_shift_reg,
	always2,
	m0_write,
	av_waitrequest_generated,
	read_latency_shift_reg_0,
	m0_write1,
	Equal22,
	always0,
	read_latency_shift_reg1,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	reset;
input 	Equal2;
input 	Equal21;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	d_read;
input 	read_accepted;
output 	read_latency_shift_reg;
input 	always2;
input 	m0_write;
output 	av_waitrequest_generated;
output 	read_latency_shift_reg_0;
input 	m0_write1;
input 	Equal22;
input 	always0;
output 	read_latency_shift_reg1;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \read_latency_shift_reg~2_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!d_read),
	.datab(!read_accepted),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \av_waitrequest_generated~0 (
	.dataa(!wait_latency_counter_0),
	.datab(!W_alu_result_4),
	.datac(!Equal2),
	.datad(!Equal21),
	.datae(!always2),
	.dataf(!m0_write),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest_generated),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest_generated~0 .extended_lut = "off";
defparam \av_waitrequest_generated~0 .lut_mask = 64'h6996966996696996;
defparam \av_waitrequest_generated~0 .shared_arith = "off";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!wait_latency_counter_0),
	.datab(!Equal22),
	.datac(!always0),
	.datad(!always2),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg1),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!wait_latency_counter_0),
	.datab(!wait_latency_counter_1),
	.datac(!always2),
	.datad(!m0_write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_0),
	.datab(!wait_latency_counter_1),
	.datac(!always2),
	.datad(!m0_write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~2 (
	.dataa(!always0),
	.datab(!read_latency_shift_reg),
	.datac(!av_waitrequest_generated),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~2 .extended_lut = "off";
defparam \read_latency_shift_reg~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \read_latency_shift_reg~2 .shared_arith = "off";

endmodule

module niosLab2_niosLab2_mm_interconnect_0_cmd_demux (
	W_alu_result_4,
	W_alu_result_3,
	Equal2,
	Equal21,
	rst1,
	av_waitrequest_generated,
	always0,
	Equal1,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	saved_grant_01,
	mem_used_11,
	WideOr0,
	Equal3,
	mem_used_12,
	av_waitrequest,
	sink_ready,
	WideOr01,
	WideOr02,
	WideOr03,
	av_waitrequest1,
	src1_valid,
	src2_valid,
	sink_ready1)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_3;
input 	Equal2;
input 	Equal21;
input 	rst1;
input 	av_waitrequest_generated;
input 	always0;
input 	Equal1;
input 	saved_grant_0;
input 	waitrequest;
input 	mem_used_1;
input 	saved_grant_01;
input 	mem_used_11;
output 	WideOr0;
input 	Equal3;
input 	mem_used_12;
input 	av_waitrequest;
output 	sink_ready;
output 	WideOr01;
output 	WideOr02;
output 	WideOr03;
input 	av_waitrequest1;
output 	src1_valid;
output 	src2_valid;
output 	sink_ready1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr0~0_combout ;
wire \WideOr0~1_combout ;


cyclonev_lcell_comb \WideOr0~2 (
	.dataa(!W_alu_result_4),
	.datab(!Equal2),
	.datac(!Equal21),
	.datad(!W_alu_result_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~2 .extended_lut = "off";
defparam \WideOr0~2 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \WideOr0~2 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~0 (
	.dataa(!Equal2),
	.datab(!Equal21),
	.datac(!Equal3),
	.datad(!mem_used_12),
	.datae(!av_waitrequest),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \sink_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~3 (
	.dataa(!Equal1),
	.datab(!\WideOr0~0_combout ),
	.datac(!\WideOr0~1_combout ),
	.datad(!WideOr0),
	.datae(!sink_ready),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr01),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~3 .extended_lut = "off";
defparam \WideOr0~3 .lut_mask = 64'hFFFFD8FFFFFFD8FF;
defparam \WideOr0~3 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~4 (
	.dataa(!Equal1),
	.datab(!\WideOr0~0_combout ),
	.datac(!\WideOr0~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr02),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~4 .extended_lut = "off";
defparam \WideOr0~4 .lut_mask = 64'h2727272727272727;
defparam \WideOr0~4 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~5 (
	.dataa(!always0),
	.datab(!av_waitrequest_generated),
	.datac(!WideOr02),
	.datad(!WideOr0),
	.datae(!sink_ready),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr03),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~5 .extended_lut = "off";
defparam \WideOr0~5 .lut_mask = 64'hFFFFFEFFFFFFFEFF;
defparam \WideOr0~5 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!W_alu_result_4),
	.datab(!Equal2),
	.datac(!Equal21),
	.datad(!W_alu_result_3),
	.datae(!av_waitrequest1),
	.dataf(!Equal1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'hFDFFFFFFFFFFFFFF;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src2_valid~0 (
	.dataa(!W_alu_result_4),
	.datab(!Equal2),
	.datac(!Equal21),
	.datad(!W_alu_result_3),
	.datae(!av_waitrequest1),
	.dataf(!Equal1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~0 .extended_lut = "off";
defparam \src2_valid~0 .lut_mask = 64'hFFFFFFFFFDFFFFFF;
defparam \src2_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~1 (
	.dataa(!Equal2),
	.datab(!Equal21),
	.datac(!Equal3),
	.datad(!av_waitrequest),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~1 .extended_lut = "off";
defparam \sink_ready~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \sink_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!saved_grant_0),
	.datab(!waitrequest),
	.datac(!mem_used_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~1 (
	.dataa(!rst1),
	.datab(!saved_grant_01),
	.datac(!mem_used_11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~1 .extended_lut = "off";
defparam \WideOr0~1 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \WideOr0~1 .shared_arith = "off";

endmodule

module niosLab2_niosLab2_mm_interconnect_0_cmd_demux_001 (
	rst1,
	i_read,
	read_accepted,
	Equal1,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	rst1;
input 	i_read;
input 	read_accepted;
input 	Equal1;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!rst1),
	.datab(!i_read),
	.datac(!read_accepted),
	.datad(!Equal1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!rst1),
	.datab(!i_read),
	.datac(!read_accepted),
	.datad(!Equal1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \src1_valid~0 .shared_arith = "off";

endmodule

module niosLab2_niosLab2_mm_interconnect_0_cmd_demux_001_1 (
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_74_0),
	.datac(!mem_56_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_74_0),
	.datac(!mem_56_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src1_valid~0 .shared_arith = "off";

endmodule

module niosLab2_niosLab2_mm_interconnect_0_cmd_demux_001_2 (
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_74_0),
	.datac(!mem_56_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_74_0),
	.datac(!mem_56_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src1_valid~0 .shared_arith = "off";

endmodule

module niosLab2_niosLab2_mm_interconnect_0_cmd_mux_001 (
	W_alu_result_4,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_7,
	W_alu_result_6,
	W_alu_result_5,
	W_alu_result_3,
	W_alu_result_2,
	F_pc_2,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_5,
	F_pc_4,
	F_pc_3,
	F_pc_1,
	F_pc_0,
	d_writedata_22,
	d_writedata_23,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_8,
	d_writedata_10,
	d_writedata_17,
	d_writedata_9,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_0,
	r_sync_rst,
	rst1,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	saved_grant_0,
	src1_valid,
	i_read,
	read_accepted,
	Equal1,
	src0_valid,
	write,
	saved_grant_1,
	src_valid,
	hbreak_enabled,
	src_data_46,
	d_byteenable_0,
	d_byteenable_2,
	d_writedata_24,
	d_byteenable_3,
	d_writedata_25,
	d_writedata_26,
	d_byteenable_1,
	d_writedata_6,
	d_writedata_7,
	src_payload,
	src_data_38,
	src_data_41,
	src_data_45,
	src_data_44,
	src_data_43,
	src_data_42,
	src_data_40,
	src_data_39,
	src_payload1,
	src_data_32,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_data_34,
	src_payload6,
	src_payload7,
	src_data_35,
	src_payload8,
	src_payload9,
	src_payload10,
	src_data_33,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_7;
input 	W_alu_result_6;
input 	W_alu_result_5;
input 	W_alu_result_3;
input 	W_alu_result_2;
input 	F_pc_2;
input 	F_pc_8;
input 	F_pc_7;
input 	F_pc_6;
input 	F_pc_5;
input 	F_pc_4;
input 	F_pc_3;
input 	F_pc_1;
input 	F_pc_0;
input 	d_writedata_22;
input 	d_writedata_23;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_16;
input 	d_writedata_8;
input 	d_writedata_10;
input 	d_writedata_17;
input 	d_writedata_9;
input 	d_writedata_18;
input 	d_writedata_19;
input 	d_writedata_20;
input 	d_writedata_21;
input 	d_writedata_0;
input 	r_sync_rst;
input 	rst1;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
output 	saved_grant_0;
input 	src1_valid;
input 	i_read;
input 	read_accepted;
input 	Equal1;
input 	src0_valid;
input 	write;
output 	saved_grant_1;
output 	src_valid;
input 	hbreak_enabled;
output 	src_data_46;
input 	d_byteenable_0;
input 	d_byteenable_2;
input 	d_writedata_24;
input 	d_byteenable_3;
input 	d_writedata_25;
input 	d_writedata_26;
input 	d_byteenable_1;
input 	d_writedata_6;
input 	d_writedata_7;
output 	src_payload;
output 	src_data_38;
output 	src_data_41;
output 	src_data_45;
output 	src_data_44;
output 	src_data_43;
output 	src_data_42;
output 	src_data_40;
output 	src_data_39;
output 	src_payload1;
output 	src_data_32;
input 	d_writedata_27;
input 	d_writedata_28;
input 	d_writedata_29;
input 	d_writedata_30;
input 	d_writedata_31;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_data_34;
output 	src_payload6;
output 	src_payload7;
output 	src_data_35;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_data_33;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


niosLab2_altera_merlin_arbitrator arb(
	.reset(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.src1_valid(src1_valid),
	.src0_valid(src0_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.write(write),
	.packet_in_progress(\packet_in_progress~q ),
	.saved_grant_1(saved_grant_1),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!rst1),
	.datab(!i_read),
	.datac(!read_accepted),
	.datad(!Equal1),
	.datae(!saved_grant_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[46] (
	.dataa(!W_alu_result_10),
	.datab(!saved_grant_0),
	.datac(!F_pc_8),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_46),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[46] .extended_lut = "off";
defparam \src_data[46] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[46] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!d_writedata_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7777777777777777;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[38] (
	.dataa(!W_alu_result_2),
	.datab(!saved_grant_0),
	.datac(!F_pc_0),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[38] .extended_lut = "off";
defparam \src_data[38] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[38] .shared_arith = "off";

cyclonev_lcell_comb \src_data[41] (
	.dataa(!W_alu_result_5),
	.datab(!saved_grant_0),
	.datac(!F_pc_3),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[41] .extended_lut = "off";
defparam \src_data[41] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[41] .shared_arith = "off";

cyclonev_lcell_comb \src_data[45] (
	.dataa(!W_alu_result_9),
	.datab(!saved_grant_0),
	.datac(!F_pc_7),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_45),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[45] .extended_lut = "off";
defparam \src_data[45] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[45] .shared_arith = "off";

cyclonev_lcell_comb \src_data[44] (
	.dataa(!W_alu_result_8),
	.datab(!saved_grant_0),
	.datac(!F_pc_6),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_44),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[44] .extended_lut = "off";
defparam \src_data[44] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[44] .shared_arith = "off";

cyclonev_lcell_comb \src_data[43] (
	.dataa(!W_alu_result_7),
	.datab(!saved_grant_0),
	.datac(!F_pc_5),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_43),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[43] .extended_lut = "off";
defparam \src_data[43] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[43] .shared_arith = "off";

cyclonev_lcell_comb \src_data[42] (
	.dataa(!W_alu_result_6),
	.datab(!saved_grant_0),
	.datac(!F_pc_4),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_42),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[42] .extended_lut = "off";
defparam \src_data[42] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[42] .shared_arith = "off";

cyclonev_lcell_comb \src_data[40] (
	.dataa(!W_alu_result_4),
	.datab(!saved_grant_0),
	.datac(!F_pc_2),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_40),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[40] .extended_lut = "off";
defparam \src_data[40] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[40] .shared_arith = "off";

cyclonev_lcell_comb \src_data[39] (
	.dataa(!W_alu_result_3),
	.datab(!saved_grant_0),
	.datac(!F_pc_1),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[39] .extended_lut = "off";
defparam \src_data[39] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[39] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!saved_grant_0),
	.datab(!hbreak_enabled),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h7777777777777777;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!d_writedata_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h7777777777777777;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!d_writedata_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h7777777777777777;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!d_writedata_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h7777777777777777;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_22),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h7777777777777777;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_23),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h7777777777777777;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_24),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h7777777777777777;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_25),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h7777777777777777;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_26),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h7777777777777777;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h7777777777777777;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h7777777777777777;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h7777777777777777;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h7777777777777777;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h7777777777777777;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h7777777777777777;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!d_writedata_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h7777777777777777;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!d_writedata_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h7777777777777777;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h7777777777777777;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h7777777777777777;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h7777777777777777;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h7777777777777777;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h7777777777777777;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_19),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h7777777777777777;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_20),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h7777777777777777;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_21),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h7777777777777777;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h7777777777777777;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h7777777777777777;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_27),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h7777777777777777;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_28),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h7777777777777777;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_29),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h7777777777777777;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h7777777777777777;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~32 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~32 .extended_lut = "off";
defparam \src_payload~32 .lut_mask = 64'h7777777777777777;
defparam \src_payload~32 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!saved_grant_0),
	.datab(!write),
	.datac(!src1_valid),
	.datad(!\packet_in_progress~q ),
	.datae(!saved_grant_1),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hFFB7FFFFFF7BFFFF;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module niosLab2_altera_merlin_arbitrator (
	reset,
	saved_grant_0,
	src1_valid,
	src0_valid,
	grant_0,
	write,
	packet_in_progress,
	saved_grant_1,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_0;
input 	src1_valid;
input 	src0_valid;
output 	grant_0;
input 	write;
input 	packet_in_progress;
input 	saved_grant_1;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~q ;
wire \top_priority_reg[1]~q ;


cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!src1_valid),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!\top_priority_reg[1]~q ),
	.datad(!src0_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \grant[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[1]~1 (
	.dataa(!src1_valid),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!\top_priority_reg[1]~q ),
	.datad(!src0_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~1 .extended_lut = "off";
defparam \grant[1]~1 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \grant[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!saved_grant_0),
	.datab(!write),
	.datac(!src1_valid),
	.datad(!src0_valid),
	.datae(!packet_in_progress),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFFFF7BB7FFFFB77B;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

endmodule

module niosLab2_niosLab2_mm_interconnect_0_cmd_mux_001_1 (
	W_alu_result_4,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_7,
	W_alu_result_6,
	W_alu_result_5,
	W_alu_result_12,
	W_alu_result_13,
	W_alu_result_14,
	W_alu_result_3,
	W_alu_result_2,
	F_pc_9,
	F_pc_10,
	F_pc_11,
	F_pc_12,
	F_pc_2,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_5,
	F_pc_4,
	F_pc_3,
	F_pc_1,
	F_pc_0,
	d_writedata_22,
	d_writedata_23,
	d_writedata_11,
	d_writedata_12,
	d_writedata_13,
	d_writedata_14,
	d_writedata_15,
	d_writedata_16,
	d_writedata_8,
	d_writedata_10,
	d_writedata_17,
	d_writedata_9,
	d_writedata_18,
	d_writedata_19,
	d_writedata_20,
	d_writedata_21,
	d_writedata_0,
	r_sync_rst,
	rst1,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	saved_grant_0,
	i_read,
	read_accepted,
	Equal1,
	src2_valid,
	src1_valid,
	read_latency_shift_reg,
	saved_grant_1,
	src_valid,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	d_byteenable_0,
	src_data_32,
	src_payload1,
	d_byteenable_2,
	src_data_34,
	src_payload2,
	d_writedata_24,
	src_payload3,
	d_byteenable_3,
	src_data_35,
	d_writedata_25,
	src_payload4,
	d_writedata_26,
	src_payload5,
	src_payload6,
	d_byteenable_1,
	src_data_33,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	d_writedata_6,
	src_payload25,
	d_writedata_7,
	src_payload26,
	d_writedata_27,
	src_payload27,
	d_writedata_28,
	src_payload28,
	d_writedata_29,
	src_payload29,
	d_writedata_30,
	src_payload30,
	d_writedata_31,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_7;
input 	W_alu_result_6;
input 	W_alu_result_5;
input 	W_alu_result_12;
input 	W_alu_result_13;
input 	W_alu_result_14;
input 	W_alu_result_3;
input 	W_alu_result_2;
input 	F_pc_9;
input 	F_pc_10;
input 	F_pc_11;
input 	F_pc_12;
input 	F_pc_2;
input 	F_pc_8;
input 	F_pc_7;
input 	F_pc_6;
input 	F_pc_5;
input 	F_pc_4;
input 	F_pc_3;
input 	F_pc_1;
input 	F_pc_0;
input 	d_writedata_22;
input 	d_writedata_23;
input 	d_writedata_11;
input 	d_writedata_12;
input 	d_writedata_13;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_16;
input 	d_writedata_8;
input 	d_writedata_10;
input 	d_writedata_17;
input 	d_writedata_9;
input 	d_writedata_18;
input 	d_writedata_19;
input 	d_writedata_20;
input 	d_writedata_21;
input 	d_writedata_0;
input 	r_sync_rst;
input 	rst1;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
output 	saved_grant_0;
input 	i_read;
input 	read_accepted;
input 	Equal1;
input 	src2_valid;
input 	src1_valid;
input 	read_latency_shift_reg;
output 	saved_grant_1;
output 	src_valid;
output 	src_payload;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_46;
output 	src_data_47;
output 	src_data_48;
output 	src_data_49;
output 	src_data_50;
input 	d_byteenable_0;
output 	src_data_32;
output 	src_payload1;
input 	d_byteenable_2;
output 	src_data_34;
output 	src_payload2;
input 	d_writedata_24;
output 	src_payload3;
input 	d_byteenable_3;
output 	src_data_35;
input 	d_writedata_25;
output 	src_payload4;
input 	d_writedata_26;
output 	src_payload5;
output 	src_payload6;
input 	d_byteenable_1;
output 	src_data_33;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
input 	d_writedata_6;
output 	src_payload25;
input 	d_writedata_7;
output 	src_payload26;
input 	d_writedata_27;
output 	src_payload27;
input 	d_writedata_28;
output 	src_payload28;
input 	d_writedata_29;
output 	src_payload29;
input 	d_writedata_30;
output 	src_payload30;
input 	d_writedata_31;
output 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


niosLab2_altera_merlin_arbitrator_1 arb(
	.reset(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.src2_valid(src2_valid),
	.src1_valid(src1_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.read_latency_shift_reg(read_latency_shift_reg),
	.packet_in_progress(\packet_in_progress~q ),
	.saved_grant_1(saved_grant_1),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!rst1),
	.datab(!i_read),
	.datac(!read_accepted),
	.datad(!Equal1),
	.datae(!saved_grant_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'hFFFDFFFFFFFDFFFF;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!d_writedata_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7777777777777777;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[38] (
	.dataa(!W_alu_result_2),
	.datab(!saved_grant_0),
	.datac(!F_pc_0),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[38] .extended_lut = "off";
defparam \src_data[38] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[38] .shared_arith = "off";

cyclonev_lcell_comb \src_data[39] (
	.dataa(!W_alu_result_3),
	.datab(!saved_grant_0),
	.datac(!F_pc_1),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[39] .extended_lut = "off";
defparam \src_data[39] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[39] .shared_arith = "off";

cyclonev_lcell_comb \src_data[40] (
	.dataa(!W_alu_result_4),
	.datab(!saved_grant_0),
	.datac(!F_pc_2),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_40),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[40] .extended_lut = "off";
defparam \src_data[40] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[40] .shared_arith = "off";

cyclonev_lcell_comb \src_data[41] (
	.dataa(!W_alu_result_5),
	.datab(!saved_grant_0),
	.datac(!F_pc_3),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[41] .extended_lut = "off";
defparam \src_data[41] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[41] .shared_arith = "off";

cyclonev_lcell_comb \src_data[42] (
	.dataa(!W_alu_result_6),
	.datab(!saved_grant_0),
	.datac(!F_pc_4),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_42),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[42] .extended_lut = "off";
defparam \src_data[42] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[42] .shared_arith = "off";

cyclonev_lcell_comb \src_data[43] (
	.dataa(!W_alu_result_7),
	.datab(!saved_grant_0),
	.datac(!F_pc_5),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_43),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[43] .extended_lut = "off";
defparam \src_data[43] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[43] .shared_arith = "off";

cyclonev_lcell_comb \src_data[44] (
	.dataa(!W_alu_result_8),
	.datab(!saved_grant_0),
	.datac(!F_pc_6),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_44),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[44] .extended_lut = "off";
defparam \src_data[44] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[44] .shared_arith = "off";

cyclonev_lcell_comb \src_data[45] (
	.dataa(!W_alu_result_9),
	.datab(!saved_grant_0),
	.datac(!F_pc_7),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_45),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[45] .extended_lut = "off";
defparam \src_data[45] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[45] .shared_arith = "off";

cyclonev_lcell_comb \src_data[46] (
	.dataa(!W_alu_result_10),
	.datab(!saved_grant_0),
	.datac(!F_pc_8),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_46),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[46] .extended_lut = "off";
defparam \src_data[46] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[46] .shared_arith = "off";

cyclonev_lcell_comb \src_data[47] (
	.dataa(!W_alu_result_11),
	.datab(!saved_grant_0),
	.datac(!F_pc_9),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_47),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[47] .extended_lut = "off";
defparam \src_data[47] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[47] .shared_arith = "off";

cyclonev_lcell_comb \src_data[48] (
	.dataa(!W_alu_result_12),
	.datab(!saved_grant_0),
	.datac(!F_pc_10),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_48),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[48] .extended_lut = "off";
defparam \src_data[48] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[48] .shared_arith = "off";

cyclonev_lcell_comb \src_data[49] (
	.dataa(!W_alu_result_13),
	.datab(!saved_grant_0),
	.datac(!F_pc_11),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_49),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[49] .extended_lut = "off";
defparam \src_data[49] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[49] .shared_arith = "off";

cyclonev_lcell_comb \src_data[50] (
	.dataa(!W_alu_result_14),
	.datab(!saved_grant_0),
	.datac(!F_pc_12),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_50),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[50] .extended_lut = "off";
defparam \src_data[50] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[50] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_22),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h7777777777777777;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_23),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h7777777777777777;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_24),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h7777777777777777;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_25),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h7777777777777777;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_26),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h7777777777777777;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h7777777777777777;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h7777777777777777;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h7777777777777777;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h7777777777777777;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h7777777777777777;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h7777777777777777;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!d_writedata_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h7777777777777777;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!d_writedata_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h7777777777777777;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!d_writedata_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h7777777777777777;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!d_writedata_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h7777777777777777;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!d_writedata_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h7777777777777777;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h7777777777777777;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h7777777777777777;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h7777777777777777;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h7777777777777777;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h7777777777777777;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_19),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h7777777777777777;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_20),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h7777777777777777;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_21),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h7777777777777777;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h7777777777777777;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h7777777777777777;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_27),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h7777777777777777;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_28),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h7777777777777777;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_29),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h7777777777777777;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h7777777777777777;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h7777777777777777;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!saved_grant_0),
	.datab(!read_latency_shift_reg),
	.datac(!src2_valid),
	.datad(!src1_valid),
	.datae(!\packet_in_progress~q ),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hFFFF7BB7FFFFB77B;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module niosLab2_altera_merlin_arbitrator_1 (
	reset,
	saved_grant_0,
	src2_valid,
	src1_valid,
	grant_0,
	read_latency_shift_reg,
	packet_in_progress,
	saved_grant_1,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_0;
input 	src2_valid;
input 	src1_valid;
output 	grant_0;
input 	read_latency_shift_reg;
input 	packet_in_progress;
input 	saved_grant_1;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~q ;
wire \top_priority_reg[1]~q ;


cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!src2_valid),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!\top_priority_reg[1]~q ),
	.datad(!src1_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \grant[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[1]~1 (
	.dataa(!src2_valid),
	.datab(!\top_priority_reg[0]~q ),
	.datac(!\top_priority_reg[1]~q ),
	.datad(!src1_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~1 .extended_lut = "off";
defparam \grant[1]~1 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \grant[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!saved_grant_0),
	.datab(!read_latency_shift_reg),
	.datac(!src2_valid),
	.datad(!src1_valid),
	.datae(!packet_in_progress),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFFFF7BB7FFFFB77B;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

endmodule

module niosLab2_niosLab2_mm_interconnect_0_router (
	W_alu_result_4,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_7,
	W_alu_result_6,
	W_alu_result_5,
	W_alu_result_12,
	W_alu_result_13,
	W_alu_result_14,
	W_alu_result_15,
	W_alu_result_16,
	W_alu_result_3,
	Equal2,
	Equal21,
	Equal22,
	Equal1,
	Equal3)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_7;
input 	W_alu_result_6;
input 	W_alu_result_5;
input 	W_alu_result_12;
input 	W_alu_result_13;
input 	W_alu_result_14;
input 	W_alu_result_15;
input 	W_alu_result_16;
input 	W_alu_result_3;
output 	Equal2;
output 	Equal21;
output 	Equal22;
output 	Equal1;
output 	Equal3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \Equal2~0 (
	.dataa(!W_alu_result_11),
	.datab(!W_alu_result_10),
	.datac(!W_alu_result_9),
	.datad(!W_alu_result_8),
	.datae(!W_alu_result_7),
	.dataf(!W_alu_result_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal2~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~1 (
	.dataa(!W_alu_result_5),
	.datab(!W_alu_result_12),
	.datac(!W_alu_result_13),
	.datad(!W_alu_result_14),
	.datae(!W_alu_result_15),
	.dataf(!W_alu_result_16),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal21),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~1 .extended_lut = "off";
defparam \Equal2~1 .lut_mask = 64'hFFFFFFFBFFFFFFFF;
defparam \Equal2~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~2 (
	.dataa(!W_alu_result_4),
	.datab(!Equal2),
	.datac(!Equal21),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal22),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~2 .extended_lut = "off";
defparam \Equal2~2 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \Equal2~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~0 (
	.dataa(!W_alu_result_11),
	.datab(!W_alu_result_12),
	.datac(!W_alu_result_13),
	.datad(!W_alu_result_14),
	.datae(!W_alu_result_15),
	.dataf(!W_alu_result_16),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hFFFFFFFDFFFFFFFF;
defparam \Equal1~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~0 (
	.dataa(!W_alu_result_4),
	.datab(!W_alu_result_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~0 .extended_lut = "off";
defparam \Equal3~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \Equal3~0 .shared_arith = "off";

endmodule

module niosLab2_niosLab2_mm_interconnect_0_router_001 (
	F_pc_9,
	F_pc_10,
	F_pc_11,
	F_pc_12,
	F_pc_14,
	F_pc_13,
	Equal1)/* synthesis synthesis_greybox=1 */;
input 	F_pc_9;
input 	F_pc_10;
input 	F_pc_11;
input 	F_pc_12;
input 	F_pc_14;
input 	F_pc_13;
output 	Equal1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \Equal1~0 (
	.dataa(!F_pc_9),
	.datab(!F_pc_10),
	.datac(!F_pc_11),
	.datad(!F_pc_12),
	.datae(!F_pc_13),
	.dataf(!F_pc_14),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hFFFDFFFFFFFFFFFF;
defparam \Equal1~0 .shared_arith = "off";

endmodule

module niosLab2_niosLab2_mm_interconnect_0_rsp_mux (
	q_a_0,
	av_readdata_pre_0,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	q_a_27,
	q_a_28,
	q_a_29,
	q_a_30,
	q_a_31,
	av_readdata_pre_7,
	av_readdata_pre_6,
	read_latency_shift_reg_0,
	src0_valid,
	read_latency_shift_reg_01,
	read_latency_shift_reg_02,
	mem_74_0,
	mem_56_0,
	WideOr1,
	src0_valid1,
	av_readdata_pre_01,
	av_readdata_pre_02,
	src_data_0,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	av_readdata_pre_11,
	av_readdata_pre_21,
	av_readdata_pre_31,
	av_readdata_pre_41,
	av_readdata_pre_51,
	av_readdata_pre_61,
	av_readdata_pre_71,
	av_readdata_pre_12,
	src_data_1,
	av_readdata_pre_22,
	src_data_2,
	av_readdata_pre_32,
	src_data_3,
	av_readdata_pre_42,
	src_data_4,
	av_readdata_pre_52,
	src_data_5,
	av_readdata_pre_27,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_30,
	av_readdata_pre_311,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9)/* synthesis synthesis_greybox=1 */;
input 	q_a_0;
input 	av_readdata_pre_0;
input 	q_a_24;
input 	q_a_25;
input 	q_a_26;
input 	q_a_1;
input 	q_a_2;
input 	q_a_3;
input 	q_a_4;
input 	q_a_5;
input 	q_a_6;
input 	q_a_7;
input 	av_readdata_pre_1;
input 	av_readdata_pre_2;
input 	av_readdata_pre_3;
input 	av_readdata_pre_4;
input 	av_readdata_pre_5;
input 	q_a_27;
input 	q_a_28;
input 	q_a_29;
input 	q_a_30;
input 	q_a_31;
input 	av_readdata_pre_7;
input 	av_readdata_pre_6;
input 	read_latency_shift_reg_0;
input 	src0_valid;
input 	read_latency_shift_reg_01;
input 	read_latency_shift_reg_02;
input 	mem_74_0;
input 	mem_56_0;
output 	WideOr1;
input 	src0_valid1;
input 	av_readdata_pre_01;
input 	av_readdata_pre_02;
output 	src_data_0;
input 	av_readdata_pre_24;
input 	av_readdata_pre_25;
input 	av_readdata_pre_26;
input 	av_readdata_pre_11;
input 	av_readdata_pre_21;
input 	av_readdata_pre_31;
input 	av_readdata_pre_41;
input 	av_readdata_pre_51;
input 	av_readdata_pre_61;
input 	av_readdata_pre_71;
input 	av_readdata_pre_12;
output 	src_data_1;
input 	av_readdata_pre_22;
output 	src_data_2;
input 	av_readdata_pre_32;
output 	src_data_3;
input 	av_readdata_pre_42;
output 	src_data_4;
input 	av_readdata_pre_52;
output 	src_data_5;
input 	av_readdata_pre_27;
input 	av_readdata_pre_28;
input 	av_readdata_pre_29;
input 	av_readdata_pre_30;
input 	av_readdata_pre_311;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \src_data[0]~0_combout ;
wire \src_data[1]~1_combout ;
wire \src_data[2]~2_combout ;
wire \src_data[3]~3_combout ;
wire \src_data[4]~4_combout ;
wire \src_data[5]~5_combout ;


cyclonev_lcell_comb \WideOr1~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!read_latency_shift_reg_01),
	.datac(!read_latency_shift_reg_02),
	.datad(!mem_74_0),
	.datae(!mem_56_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr1),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr1~0 .extended_lut = "off";
defparam \WideOr1~0 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \WideOr1~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0] (
	.dataa(!src0_valid1),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_01),
	.datad(!q_a_0),
	.datae(!\src_data[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0] .extended_lut = "off";
defparam \src_data[0] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[0] .shared_arith = "off";

cyclonev_lcell_comb \src_data[1] (
	.dataa(!src0_valid1),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_11),
	.datad(!q_a_1),
	.datae(!\src_data[1]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1] .extended_lut = "off";
defparam \src_data[1] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[1] .shared_arith = "off";

cyclonev_lcell_comb \src_data[2] (
	.dataa(!src0_valid1),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_21),
	.datad(!q_a_2),
	.datae(!\src_data[2]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2] .extended_lut = "off";
defparam \src_data[2] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[2] .shared_arith = "off";

cyclonev_lcell_comb \src_data[3] (
	.dataa(!src0_valid1),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_31),
	.datad(!q_a_3),
	.datae(!\src_data[3]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3] .extended_lut = "off";
defparam \src_data[3] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[3] .shared_arith = "off";

cyclonev_lcell_comb \src_data[4] (
	.dataa(!src0_valid1),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_41),
	.datad(!q_a_4),
	.datae(!\src_data[4]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4] .extended_lut = "off";
defparam \src_data[4] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[4] .shared_arith = "off";

cyclonev_lcell_comb \src_data[5] (
	.dataa(!src0_valid1),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_51),
	.datad(!q_a_5),
	.datae(!\src_data[5]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5] .extended_lut = "off";
defparam \src_data[5] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[5] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid1),
	.datac(!src0_valid),
	.datad(!av_readdata_pre_71),
	.datae(!q_a_7),
	.dataf(!av_readdata_pre_7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid1),
	.datac(!src0_valid),
	.datad(!av_readdata_pre_61),
	.datae(!q_a_6),
	.dataf(!av_readdata_pre_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!src0_valid1),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_24),
	.datad(!q_a_24),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!src0_valid1),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_25),
	.datad(!q_a_25),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!src0_valid1),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_27),
	.datad(!q_a_27),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!src0_valid1),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_26),
	.datad(!q_a_26),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!src0_valid1),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_311),
	.datad(!q_a_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!src0_valid1),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_30),
	.datad(!q_a_30),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!src0_valid1),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_28),
	.datad(!q_a_28),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!src0_valid1),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_29),
	.datad(!q_a_29),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!read_latency_shift_reg_01),
	.datac(!av_readdata_pre_0),
	.datad(!av_readdata_pre_02),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~0 .extended_lut = "off";
defparam \src_data[0]~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!read_latency_shift_reg_01),
	.datac(!av_readdata_pre_1),
	.datad(!av_readdata_pre_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~1 .extended_lut = "off";
defparam \src_data[1]~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~2 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!read_latency_shift_reg_01),
	.datac(!av_readdata_pre_2),
	.datad(!av_readdata_pre_22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~2 .extended_lut = "off";
defparam \src_data[2]~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~3 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!read_latency_shift_reg_01),
	.datac(!av_readdata_pre_3),
	.datad(!av_readdata_pre_32),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~3 .extended_lut = "off";
defparam \src_data[3]~3 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4]~4 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!read_latency_shift_reg_01),
	.datac(!av_readdata_pre_4),
	.datad(!av_readdata_pre_42),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4]~4 .extended_lut = "off";
defparam \src_data[4]~4 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~5 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!read_latency_shift_reg_01),
	.datac(!av_readdata_pre_5),
	.datad(!av_readdata_pre_52),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~5 .extended_lut = "off";
defparam \src_data[5]~5 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[5]~5 .shared_arith = "off";

endmodule

module niosLab2_niosLab2_mm_interconnect_0_rsp_mux_001 (
	q_a_0,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_12,
	q_a_14,
	q_a_2,
	q_a_8,
	q_a_10,
	q_a_17,
	q_a_9,
	q_a_6,
	q_a_7,
	q_a_27,
	q_a_28,
	q_a_29,
	q_a_30,
	q_a_31,
	av_readdata_pre_0,
	av_readdata_pre_22,
	src1_valid,
	src1_valid1,
	src_data_22,
	av_readdata_pre_23,
	src_data_23,
	av_readdata_pre_24,
	src_data_24,
	av_readdata_pre_25,
	src_data_25,
	av_readdata_pre_26,
	src_data_26,
	av_readdata_pre_12,
	src_data_12,
	av_readdata_pre_14,
	src_data_14,
	src_data_0,
	av_readdata_pre_2,
	src_data_2,
	av_readdata_pre_8,
	src_data_8,
	av_readdata_pre_10,
	src_data_10,
	av_readdata_pre_17,
	src_data_17,
	av_readdata_pre_9,
	src_data_9,
	av_readdata_pre_6,
	src_data_6,
	av_readdata_pre_7,
	src_data_7,
	av_readdata_pre_27,
	src_data_27,
	av_readdata_pre_28,
	src_data_28,
	av_readdata_pre_29,
	src_data_29,
	av_readdata_pre_30,
	src_data_30,
	av_readdata_pre_31,
	src_data_31)/* synthesis synthesis_greybox=1 */;
input 	q_a_0;
input 	q_a_22;
input 	q_a_23;
input 	q_a_24;
input 	q_a_25;
input 	q_a_26;
input 	q_a_12;
input 	q_a_14;
input 	q_a_2;
input 	q_a_8;
input 	q_a_10;
input 	q_a_17;
input 	q_a_9;
input 	q_a_6;
input 	q_a_7;
input 	q_a_27;
input 	q_a_28;
input 	q_a_29;
input 	q_a_30;
input 	q_a_31;
input 	av_readdata_pre_0;
input 	av_readdata_pre_22;
input 	src1_valid;
input 	src1_valid1;
output 	src_data_22;
input 	av_readdata_pre_23;
output 	src_data_23;
input 	av_readdata_pre_24;
output 	src_data_24;
input 	av_readdata_pre_25;
output 	src_data_25;
input 	av_readdata_pre_26;
output 	src_data_26;
input 	av_readdata_pre_12;
output 	src_data_12;
input 	av_readdata_pre_14;
output 	src_data_14;
output 	src_data_0;
input 	av_readdata_pre_2;
output 	src_data_2;
input 	av_readdata_pre_8;
output 	src_data_8;
input 	av_readdata_pre_10;
output 	src_data_10;
input 	av_readdata_pre_17;
output 	src_data_17;
input 	av_readdata_pre_9;
output 	src_data_9;
input 	av_readdata_pre_6;
output 	src_data_6;
input 	av_readdata_pre_7;
output 	src_data_7;
input 	av_readdata_pre_27;
output 	src_data_27;
input 	av_readdata_pre_28;
output 	src_data_28;
input 	av_readdata_pre_29;
output 	src_data_29;
input 	av_readdata_pre_30;
output 	src_data_30;
input 	av_readdata_pre_31;
output 	src_data_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src_data[22] (
	.dataa(!av_readdata_pre_22),
	.datab(!src1_valid),
	.datac(!q_a_22),
	.datad(!src1_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[22] .extended_lut = "off";
defparam \src_data[22] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[22] .shared_arith = "off";

cyclonev_lcell_comb \src_data[23] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_23),
	.datad(!q_a_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[23] .extended_lut = "off";
defparam \src_data[23] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[23] .shared_arith = "off";

cyclonev_lcell_comb \src_data[24] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_24),
	.datad(!q_a_24),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[24] .extended_lut = "off";
defparam \src_data[24] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[24] .shared_arith = "off";

cyclonev_lcell_comb \src_data[25] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_25),
	.datad(!q_a_25),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[25] .extended_lut = "off";
defparam \src_data[25] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[25] .shared_arith = "off";

cyclonev_lcell_comb \src_data[26] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_26),
	.datad(!q_a_26),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[26] .extended_lut = "off";
defparam \src_data[26] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[26] .shared_arith = "off";

cyclonev_lcell_comb \src_data[12] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_12),
	.datad(!q_a_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[12] .extended_lut = "off";
defparam \src_data[12] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[12] .shared_arith = "off";

cyclonev_lcell_comb \src_data[14] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_14),
	.datad(!q_a_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[14] .extended_lut = "off";
defparam \src_data[14] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[14] .shared_arith = "off";

cyclonev_lcell_comb \src_data[0] (
	.dataa(!av_readdata_pre_0),
	.datab(!q_a_0),
	.datac(!src1_valid),
	.datad(!src1_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0] .extended_lut = "off";
defparam \src_data[0] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[0] .shared_arith = "off";

cyclonev_lcell_comb \src_data[2] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_2),
	.datad(!q_a_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2] .extended_lut = "off";
defparam \src_data[2] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[2] .shared_arith = "off";

cyclonev_lcell_comb \src_data[8] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_8),
	.datad(!q_a_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8] .extended_lut = "off";
defparam \src_data[8] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[8] .shared_arith = "off";

cyclonev_lcell_comb \src_data[10] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_10),
	.datad(!q_a_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[10] .extended_lut = "off";
defparam \src_data[10] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[10] .shared_arith = "off";

cyclonev_lcell_comb \src_data[17] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_17),
	.datad(!q_a_17),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[17] .extended_lut = "off";
defparam \src_data[17] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[17] .shared_arith = "off";

cyclonev_lcell_comb \src_data[9] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_9),
	.datad(!q_a_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9] .extended_lut = "off";
defparam \src_data[9] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[9] .shared_arith = "off";

cyclonev_lcell_comb \src_data[6] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_6),
	.datad(!q_a_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6] .extended_lut = "off";
defparam \src_data[6] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[6] .shared_arith = "off";

cyclonev_lcell_comb \src_data[7] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_7),
	.datad(!q_a_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7] .extended_lut = "off";
defparam \src_data[7] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[7] .shared_arith = "off";

cyclonev_lcell_comb \src_data[27] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_27),
	.datad(!q_a_27),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[27] .extended_lut = "off";
defparam \src_data[27] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[27] .shared_arith = "off";

cyclonev_lcell_comb \src_data[28] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_28),
	.datad(!q_a_28),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[28] .extended_lut = "off";
defparam \src_data[28] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[28] .shared_arith = "off";

cyclonev_lcell_comb \src_data[29] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_29),
	.datad(!q_a_29),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[29] .extended_lut = "off";
defparam \src_data[29] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[29] .shared_arith = "off";

cyclonev_lcell_comb \src_data[30] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_30),
	.datad(!q_a_30),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[30] .extended_lut = "off";
defparam \src_data[30] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[30] .shared_arith = "off";

cyclonev_lcell_comb \src_data[31] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_31),
	.datad(!q_a_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[31] .extended_lut = "off";
defparam \src_data[31] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[31] .shared_arith = "off";

endmodule

module niosLab2_niosLab2_nios2_gen2_0 (
	W_alu_result_4,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_7,
	W_alu_result_6,
	W_alu_result_5,
	W_alu_result_12,
	W_alu_result_13,
	W_alu_result_14,
	W_alu_result_15,
	W_alu_result_16,
	W_alu_result_3,
	W_alu_result_2,
	F_pc_9,
	F_pc_10,
	F_pc_11,
	F_pc_12,
	F_pc_14,
	q_a_22,
	q_a_23,
	q_a_11,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_15,
	q_a_16,
	q_a_1,
	q_a_3,
	q_a_4,
	q_a_5,
	F_pc_2,
	q_a_8,
	q_a_10,
	q_a_17,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_5,
	F_pc_4,
	F_pc_3,
	q_a_9,
	q_a_18,
	q_a_19,
	q_a_20,
	q_a_21,
	F_pc_1,
	F_pc_0,
	readdata_0,
	readdata_22,
	d_writedata_22,
	readdata_23,
	d_writedata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_11,
	d_writedata_11,
	readdata_12,
	d_writedata_12,
	readdata_13,
	d_writedata_13,
	readdata_14,
	d_writedata_14,
	readdata_15,
	d_writedata_15,
	readdata_16,
	d_writedata_16,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_8,
	d_writedata_8,
	readdata_10,
	d_writedata_10,
	readdata_17,
	d_writedata_17,
	readdata_9,
	d_writedata_9,
	readdata_18,
	d_writedata_18,
	readdata_19,
	d_writedata_19,
	readdata_20,
	d_writedata_20,
	readdata_21,
	d_writedata_21,
	av_readdata_pre_16,
	readdata_6,
	readdata_7,
	readdata_27,
	readdata_28,
	readdata_29,
	readdata_30,
	readdata_31,
	av_readdata_pre_19,
	av_readdata_pre_18,
	av_readdata_pre_17,
	av_readdata_pre_20,
	av_readdata_pre_21,
	av_readdata_pre_22,
	av_waitrequest,
	sr_0,
	ir_out_0,
	ir_out_1,
	d_writedata_0,
	r_sync_rst,
	d_write,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_read,
	always2,
	av_waitrequest1,
	read_latency_shift_reg,
	saved_grant_0,
	debug_mem_slave_waitrequest,
	mem_used_1,
	WideOr0,
	src0_valid,
	read_latency_shift_reg_0,
	WideOr1,
	src1_valid,
	i_read,
	F_pc_13,
	src_valid,
	mem,
	hbreak_enabled,
	av_waitrequest2,
	src0_valid1,
	src_data_0,
	av_readdata_pre_221,
	src1_valid1,
	src1_valid2,
	src_data_22,
	av_readdata_pre_23,
	src_data_23,
	src_data_24,
	src_data_25,
	src_data_26,
	av_readdata_pre_11,
	av_readdata_pre_12,
	src_data_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	src_data_14,
	av_readdata_pre_15,
	av_readdata_pre_161,
	src_data_01,
	av_readdata_pre_1,
	src_data_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_8,
	src_data_8,
	av_readdata_pre_10,
	src_data_10,
	av_readdata_pre_171,
	src_data_17,
	av_readdata_pre_9,
	src_data_9,
	av_readdata_pre_181,
	av_readdata_pre_191,
	av_readdata_pre_201,
	av_readdata_pre_211,
	src_data_6,
	src_data_46,
	src_data_7,
	src_data_1,
	src_data_21,
	src_data_3,
	src_data_4,
	src_data_5,
	r_early_rst,
	d_byteenable_0,
	av_readdata_pre_81,
	d_byteenable_2,
	d_writedata_24,
	d_byteenable_3,
	d_writedata_25,
	d_writedata_26,
	d_byteenable_1,
	src_data_27,
	src_data_28,
	src_data_29,
	src_data_30,
	src_data_31,
	av_readdata_pre_101,
	av_readdata_pre_91,
	src_payload,
	src_payload1,
	av_readdata_pre_121,
	av_readdata_pre_131,
	av_readdata_pre_141,
	av_readdata_pre_151,
	d_writedata_6,
	d_writedata_7,
	src_payload2,
	src_data_38,
	src_data_41,
	src_data_45,
	src_data_44,
	src_data_43,
	src_data_42,
	src_data_40,
	src_data_39,
	src_payload3,
	src_data_32,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_data_34,
	src_payload16,
	src_payload17,
	src_data_35,
	src_payload18,
	src_payload19,
	src_payload20,
	src_data_33,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_payload41,
	src_payload42,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	W_alu_result_4;
output 	W_alu_result_11;
output 	W_alu_result_10;
output 	W_alu_result_9;
output 	W_alu_result_8;
output 	W_alu_result_7;
output 	W_alu_result_6;
output 	W_alu_result_5;
output 	W_alu_result_12;
output 	W_alu_result_13;
output 	W_alu_result_14;
output 	W_alu_result_15;
output 	W_alu_result_16;
output 	W_alu_result_3;
output 	W_alu_result_2;
output 	F_pc_9;
output 	F_pc_10;
output 	F_pc_11;
output 	F_pc_12;
output 	F_pc_14;
input 	q_a_22;
input 	q_a_23;
input 	q_a_11;
input 	q_a_12;
input 	q_a_13;
input 	q_a_14;
input 	q_a_15;
input 	q_a_16;
input 	q_a_1;
input 	q_a_3;
input 	q_a_4;
input 	q_a_5;
output 	F_pc_2;
input 	q_a_8;
input 	q_a_10;
input 	q_a_17;
output 	F_pc_8;
output 	F_pc_7;
output 	F_pc_6;
output 	F_pc_5;
output 	F_pc_4;
output 	F_pc_3;
input 	q_a_9;
input 	q_a_18;
input 	q_a_19;
input 	q_a_20;
input 	q_a_21;
output 	F_pc_1;
output 	F_pc_0;
output 	readdata_0;
output 	readdata_22;
output 	d_writedata_22;
output 	readdata_23;
output 	d_writedata_23;
output 	readdata_24;
output 	readdata_25;
output 	readdata_26;
output 	readdata_11;
output 	d_writedata_11;
output 	readdata_12;
output 	d_writedata_12;
output 	readdata_13;
output 	d_writedata_13;
output 	readdata_14;
output 	d_writedata_14;
output 	readdata_15;
output 	d_writedata_15;
output 	readdata_16;
output 	d_writedata_16;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_8;
output 	d_writedata_8;
output 	readdata_10;
output 	d_writedata_10;
output 	readdata_17;
output 	d_writedata_17;
output 	readdata_9;
output 	d_writedata_9;
output 	readdata_18;
output 	d_writedata_18;
output 	readdata_19;
output 	d_writedata_19;
output 	readdata_20;
output 	d_writedata_20;
output 	readdata_21;
output 	d_writedata_21;
input 	av_readdata_pre_16;
output 	readdata_6;
output 	readdata_7;
output 	readdata_27;
output 	readdata_28;
output 	readdata_29;
output 	readdata_30;
output 	readdata_31;
input 	av_readdata_pre_19;
input 	av_readdata_pre_18;
input 	av_readdata_pre_17;
input 	av_readdata_pre_20;
input 	av_readdata_pre_21;
input 	av_readdata_pre_22;
input 	av_waitrequest;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
output 	d_writedata_0;
input 	r_sync_rst;
output 	d_write;
output 	d_writedata_1;
output 	d_writedata_2;
output 	d_writedata_3;
output 	d_writedata_4;
output 	d_writedata_5;
output 	d_read;
input 	always2;
input 	av_waitrequest1;
input 	read_latency_shift_reg;
input 	saved_grant_0;
output 	debug_mem_slave_waitrequest;
input 	mem_used_1;
input 	WideOr0;
input 	src0_valid;
input 	read_latency_shift_reg_0;
input 	WideOr1;
input 	src1_valid;
output 	i_read;
output 	F_pc_13;
input 	src_valid;
input 	mem;
output 	hbreak_enabled;
input 	av_waitrequest2;
input 	src0_valid1;
input 	src_data_0;
input 	av_readdata_pre_221;
input 	src1_valid1;
input 	src1_valid2;
input 	src_data_22;
input 	av_readdata_pre_23;
input 	src_data_23;
input 	src_data_24;
input 	src_data_25;
input 	src_data_26;
input 	av_readdata_pre_11;
input 	av_readdata_pre_12;
input 	src_data_12;
input 	av_readdata_pre_13;
input 	av_readdata_pre_14;
input 	src_data_14;
input 	av_readdata_pre_15;
input 	av_readdata_pre_161;
input 	src_data_01;
input 	av_readdata_pre_1;
input 	src_data_2;
input 	av_readdata_pre_3;
input 	av_readdata_pre_4;
input 	av_readdata_pre_5;
input 	av_readdata_pre_8;
input 	src_data_8;
input 	av_readdata_pre_10;
input 	src_data_10;
input 	av_readdata_pre_171;
input 	src_data_17;
input 	av_readdata_pre_9;
input 	src_data_9;
input 	av_readdata_pre_181;
input 	av_readdata_pre_191;
input 	av_readdata_pre_201;
input 	av_readdata_pre_211;
input 	src_data_6;
input 	src_data_46;
input 	src_data_7;
input 	src_data_1;
input 	src_data_21;
input 	src_data_3;
input 	src_data_4;
input 	src_data_5;
input 	r_early_rst;
output 	d_byteenable_0;
input 	av_readdata_pre_81;
output 	d_byteenable_2;
output 	d_writedata_24;
output 	d_byteenable_3;
output 	d_writedata_25;
output 	d_writedata_26;
output 	d_byteenable_1;
input 	src_data_27;
input 	src_data_28;
input 	src_data_29;
input 	src_data_30;
input 	src_data_31;
input 	av_readdata_pre_101;
input 	av_readdata_pre_91;
input 	src_payload;
input 	src_payload1;
input 	av_readdata_pre_121;
input 	av_readdata_pre_131;
input 	av_readdata_pre_141;
input 	av_readdata_pre_151;
output 	d_writedata_6;
output 	d_writedata_7;
input 	src_payload2;
input 	src_data_38;
input 	src_data_41;
input 	src_data_45;
input 	src_data_44;
input 	src_data_43;
input 	src_data_42;
input 	src_data_40;
input 	src_data_39;
input 	src_payload3;
input 	src_data_32;
output 	d_writedata_27;
output 	d_writedata_28;
output 	d_writedata_29;
output 	d_writedata_30;
output 	d_writedata_31;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_data_34;
input 	src_payload16;
input 	src_payload17;
input 	src_data_35;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_data_33;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	src_payload33;
input 	src_payload34;
input 	src_payload35;
input 	src_payload36;
input 	src_payload37;
input 	src_payload38;
input 	src_payload39;
input 	src_payload40;
input 	src_payload41;
input 	src_payload42;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosLab2_niosLab2_nios2_gen2_0_cpu cpu(
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_16(W_alu_result_16),
	.W_alu_result_3(W_alu_result_3),
	.W_alu_result_2(W_alu_result_2),
	.F_pc_9(F_pc_9),
	.F_pc_10(F_pc_10),
	.F_pc_11(F_pc_11),
	.F_pc_12(F_pc_12),
	.F_pc_14(F_pc_14),
	.q_a_22(q_a_22),
	.q_a_23(q_a_23),
	.q_a_11(q_a_11),
	.q_a_12(q_a_12),
	.q_a_13(q_a_13),
	.q_a_14(q_a_14),
	.q_a_15(q_a_15),
	.q_a_16(q_a_16),
	.q_a_1(q_a_1),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.F_pc_2(F_pc_2),
	.q_a_8(q_a_8),
	.q_a_10(q_a_10),
	.q_a_17(q_a_17),
	.F_pc_8(F_pc_8),
	.F_pc_7(F_pc_7),
	.F_pc_6(F_pc_6),
	.F_pc_5(F_pc_5),
	.F_pc_4(F_pc_4),
	.F_pc_3(F_pc_3),
	.q_a_9(q_a_9),
	.q_a_18(q_a_18),
	.q_a_19(q_a_19),
	.q_a_20(q_a_20),
	.q_a_21(q_a_21),
	.F_pc_1(F_pc_1),
	.F_pc_0(F_pc_0),
	.readdata_0(readdata_0),
	.readdata_22(readdata_22),
	.d_writedata_22(d_writedata_22),
	.readdata_23(readdata_23),
	.d_writedata_23(d_writedata_23),
	.readdata_24(readdata_24),
	.readdata_25(readdata_25),
	.readdata_26(readdata_26),
	.readdata_11(readdata_11),
	.d_writedata_11(d_writedata_11),
	.readdata_12(readdata_12),
	.d_writedata_12(d_writedata_12),
	.readdata_13(readdata_13),
	.d_writedata_13(d_writedata_13),
	.readdata_14(readdata_14),
	.d_writedata_14(d_writedata_14),
	.readdata_15(readdata_15),
	.d_writedata_15(d_writedata_15),
	.readdata_16(readdata_16),
	.d_writedata_16(d_writedata_16),
	.readdata_1(readdata_1),
	.readdata_2(readdata_2),
	.readdata_3(readdata_3),
	.readdata_4(readdata_4),
	.readdata_5(readdata_5),
	.readdata_8(readdata_8),
	.d_writedata_8(d_writedata_8),
	.readdata_10(readdata_10),
	.d_writedata_10(d_writedata_10),
	.readdata_17(readdata_17),
	.d_writedata_17(d_writedata_17),
	.readdata_9(readdata_9),
	.d_writedata_9(d_writedata_9),
	.readdata_18(readdata_18),
	.d_writedata_18(d_writedata_18),
	.readdata_19(readdata_19),
	.d_writedata_19(d_writedata_19),
	.readdata_20(readdata_20),
	.d_writedata_20(d_writedata_20),
	.readdata_21(readdata_21),
	.d_writedata_21(d_writedata_21),
	.av_readdata_pre_16(av_readdata_pre_16),
	.readdata_6(readdata_6),
	.readdata_7(readdata_7),
	.readdata_27(readdata_27),
	.readdata_28(readdata_28),
	.readdata_29(readdata_29),
	.readdata_30(readdata_30),
	.readdata_31(readdata_31),
	.av_readdata_pre_19(av_readdata_pre_19),
	.av_readdata_pre_18(av_readdata_pre_18),
	.av_readdata_pre_17(av_readdata_pre_17),
	.av_readdata_pre_20(av_readdata_pre_20),
	.av_readdata_pre_21(av_readdata_pre_21),
	.av_readdata_pre_22(av_readdata_pre_22),
	.av_waitrequest(av_waitrequest),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.d_write1(d_write),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_read1(d_read),
	.always2(always2),
	.av_waitrequest1(av_waitrequest1),
	.read_latency_shift_reg(read_latency_shift_reg),
	.saved_grant_0(saved_grant_0),
	.debug_mem_slave_waitrequest(debug_mem_slave_waitrequest),
	.mem_used_1(mem_used_1),
	.WideOr0(WideOr0),
	.src0_valid(src0_valid),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.WideOr1(WideOr1),
	.src1_valid(src1_valid),
	.i_read1(i_read),
	.F_pc_13(F_pc_13),
	.src_valid(src_valid),
	.mem(mem),
	.hbreak_enabled1(hbreak_enabled),
	.av_waitrequest2(av_waitrequest2),
	.src0_valid1(src0_valid1),
	.src_data_0(src_data_0),
	.av_readdata_pre_221(av_readdata_pre_221),
	.src1_valid1(src1_valid1),
	.src1_valid2(src1_valid2),
	.src_data_22(src_data_22),
	.av_readdata_pre_23(av_readdata_pre_23),
	.src_data_23(src_data_23),
	.src_data_24(src_data_24),
	.src_data_25(src_data_25),
	.src_data_26(src_data_26),
	.av_readdata_pre_11(av_readdata_pre_11),
	.av_readdata_pre_12(av_readdata_pre_12),
	.src_data_12(src_data_12),
	.av_readdata_pre_13(av_readdata_pre_13),
	.av_readdata_pre_14(av_readdata_pre_14),
	.src_data_14(src_data_14),
	.av_readdata_pre_15(av_readdata_pre_15),
	.av_readdata_pre_161(av_readdata_pre_161),
	.src_data_01(src_data_01),
	.av_readdata_pre_1(av_readdata_pre_1),
	.src_data_2(src_data_2),
	.av_readdata_pre_3(av_readdata_pre_3),
	.av_readdata_pre_4(av_readdata_pre_4),
	.av_readdata_pre_5(av_readdata_pre_5),
	.av_readdata_pre_8(av_readdata_pre_8),
	.src_data_8(src_data_8),
	.av_readdata_pre_10(av_readdata_pre_10),
	.src_data_10(src_data_10),
	.av_readdata_pre_171(av_readdata_pre_171),
	.src_data_17(src_data_17),
	.av_readdata_pre_9(av_readdata_pre_9),
	.src_data_9(src_data_9),
	.av_readdata_pre_181(av_readdata_pre_181),
	.av_readdata_pre_191(av_readdata_pre_191),
	.av_readdata_pre_201(av_readdata_pre_201),
	.av_readdata_pre_211(av_readdata_pre_211),
	.src_data_6(src_data_6),
	.src_data_46(src_data_46),
	.src_data_7(src_data_7),
	.src_data_1(src_data_1),
	.src_data_21(src_data_21),
	.src_data_3(src_data_3),
	.src_data_4(src_data_4),
	.src_data_5(src_data_5),
	.r_early_rst(r_early_rst),
	.d_byteenable_0(d_byteenable_0),
	.av_readdata_pre_81(av_readdata_pre_81),
	.d_byteenable_2(d_byteenable_2),
	.d_writedata_24(d_writedata_24),
	.d_byteenable_3(d_byteenable_3),
	.d_writedata_25(d_writedata_25),
	.d_writedata_26(d_writedata_26),
	.d_byteenable_1(d_byteenable_1),
	.src_data_27(src_data_27),
	.src_data_28(src_data_28),
	.src_data_29(src_data_29),
	.src_data_30(src_data_30),
	.src_data_31(src_data_31),
	.av_readdata_pre_101(av_readdata_pre_101),
	.av_readdata_pre_91(av_readdata_pre_91),
	.src_payload(src_payload),
	.src_payload1(src_payload1),
	.av_readdata_pre_121(av_readdata_pre_121),
	.av_readdata_pre_131(av_readdata_pre_131),
	.av_readdata_pre_141(av_readdata_pre_141),
	.av_readdata_pre_151(av_readdata_pre_151),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.src_payload2(src_payload2),
	.src_data_38(src_data_38),
	.src_data_41(src_data_41),
	.src_data_45(src_data_45),
	.src_data_44(src_data_44),
	.src_data_43(src_data_43),
	.src_data_42(src_data_42),
	.src_data_40(src_data_40),
	.src_data_39(src_data_39),
	.src_payload3(src_payload3),
	.src_data_32(src_data_32),
	.d_writedata_27(d_writedata_27),
	.d_writedata_28(d_writedata_28),
	.d_writedata_29(d_writedata_29),
	.d_writedata_30(d_writedata_30),
	.d_writedata_31(d_writedata_31),
	.src_payload4(src_payload4),
	.src_payload5(src_payload5),
	.src_payload6(src_payload6),
	.src_payload7(src_payload7),
	.src_payload8(src_payload8),
	.src_payload9(src_payload9),
	.src_payload10(src_payload10),
	.src_payload11(src_payload11),
	.src_payload12(src_payload12),
	.src_payload13(src_payload13),
	.src_payload14(src_payload14),
	.src_payload15(src_payload15),
	.src_data_34(src_data_34),
	.src_payload16(src_payload16),
	.src_payload17(src_payload17),
	.src_data_35(src_data_35),
	.src_payload18(src_payload18),
	.src_payload19(src_payload19),
	.src_payload20(src_payload20),
	.src_data_33(src_data_33),
	.src_payload21(src_payload21),
	.src_payload22(src_payload22),
	.src_payload23(src_payload23),
	.src_payload24(src_payload24),
	.src_payload25(src_payload25),
	.src_payload26(src_payload26),
	.src_payload27(src_payload27),
	.src_payload28(src_payload28),
	.src_payload29(src_payload29),
	.src_payload30(src_payload30),
	.src_payload31(src_payload31),
	.src_payload32(src_payload32),
	.src_payload33(src_payload33),
	.src_payload34(src_payload34),
	.src_payload35(src_payload35),
	.src_payload36(src_payload36),
	.src_payload37(src_payload37),
	.src_payload38(src_payload38),
	.src_payload39(src_payload39),
	.src_payload40(src_payload40),
	.src_payload41(src_payload41),
	.src_payload42(src_payload42),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

endmodule

module niosLab2_niosLab2_nios2_gen2_0_cpu (
	W_alu_result_4,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_7,
	W_alu_result_6,
	W_alu_result_5,
	W_alu_result_12,
	W_alu_result_13,
	W_alu_result_14,
	W_alu_result_15,
	W_alu_result_16,
	W_alu_result_3,
	W_alu_result_2,
	F_pc_9,
	F_pc_10,
	F_pc_11,
	F_pc_12,
	F_pc_14,
	q_a_22,
	q_a_23,
	q_a_11,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_15,
	q_a_16,
	q_a_1,
	q_a_3,
	q_a_4,
	q_a_5,
	F_pc_2,
	q_a_8,
	q_a_10,
	q_a_17,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_5,
	F_pc_4,
	F_pc_3,
	q_a_9,
	q_a_18,
	q_a_19,
	q_a_20,
	q_a_21,
	F_pc_1,
	F_pc_0,
	readdata_0,
	readdata_22,
	d_writedata_22,
	readdata_23,
	d_writedata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_11,
	d_writedata_11,
	readdata_12,
	d_writedata_12,
	readdata_13,
	d_writedata_13,
	readdata_14,
	d_writedata_14,
	readdata_15,
	d_writedata_15,
	readdata_16,
	d_writedata_16,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_8,
	d_writedata_8,
	readdata_10,
	d_writedata_10,
	readdata_17,
	d_writedata_17,
	readdata_9,
	d_writedata_9,
	readdata_18,
	d_writedata_18,
	readdata_19,
	d_writedata_19,
	readdata_20,
	d_writedata_20,
	readdata_21,
	d_writedata_21,
	av_readdata_pre_16,
	readdata_6,
	readdata_7,
	readdata_27,
	readdata_28,
	readdata_29,
	readdata_30,
	readdata_31,
	av_readdata_pre_19,
	av_readdata_pre_18,
	av_readdata_pre_17,
	av_readdata_pre_20,
	av_readdata_pre_21,
	av_readdata_pre_22,
	av_waitrequest,
	sr_0,
	ir_out_0,
	ir_out_1,
	d_writedata_0,
	r_sync_rst,
	d_write1,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_read1,
	always2,
	av_waitrequest1,
	read_latency_shift_reg,
	saved_grant_0,
	debug_mem_slave_waitrequest,
	mem_used_1,
	WideOr0,
	src0_valid,
	read_latency_shift_reg_0,
	WideOr1,
	src1_valid,
	i_read1,
	F_pc_13,
	src_valid,
	mem,
	hbreak_enabled1,
	av_waitrequest2,
	src0_valid1,
	src_data_0,
	av_readdata_pre_221,
	src1_valid1,
	src1_valid2,
	src_data_22,
	av_readdata_pre_23,
	src_data_23,
	src_data_24,
	src_data_25,
	src_data_26,
	av_readdata_pre_11,
	av_readdata_pre_12,
	src_data_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	src_data_14,
	av_readdata_pre_15,
	av_readdata_pre_161,
	src_data_01,
	av_readdata_pre_1,
	src_data_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_8,
	src_data_8,
	av_readdata_pre_10,
	src_data_10,
	av_readdata_pre_171,
	src_data_17,
	av_readdata_pre_9,
	src_data_9,
	av_readdata_pre_181,
	av_readdata_pre_191,
	av_readdata_pre_201,
	av_readdata_pre_211,
	src_data_6,
	src_data_46,
	src_data_7,
	src_data_1,
	src_data_21,
	src_data_3,
	src_data_4,
	src_data_5,
	r_early_rst,
	d_byteenable_0,
	av_readdata_pre_81,
	d_byteenable_2,
	d_writedata_24,
	d_byteenable_3,
	d_writedata_25,
	d_writedata_26,
	d_byteenable_1,
	src_data_27,
	src_data_28,
	src_data_29,
	src_data_30,
	src_data_31,
	av_readdata_pre_101,
	av_readdata_pre_91,
	src_payload,
	src_payload1,
	av_readdata_pre_121,
	av_readdata_pre_131,
	av_readdata_pre_141,
	av_readdata_pre_151,
	d_writedata_6,
	d_writedata_7,
	src_payload2,
	src_data_38,
	src_data_41,
	src_data_45,
	src_data_44,
	src_data_43,
	src_data_42,
	src_data_40,
	src_data_39,
	src_payload3,
	src_data_32,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_data_34,
	src_payload16,
	src_payload17,
	src_data_35,
	src_payload18,
	src_payload19,
	src_payload20,
	src_data_33,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_payload41,
	src_payload42,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	W_alu_result_4;
output 	W_alu_result_11;
output 	W_alu_result_10;
output 	W_alu_result_9;
output 	W_alu_result_8;
output 	W_alu_result_7;
output 	W_alu_result_6;
output 	W_alu_result_5;
output 	W_alu_result_12;
output 	W_alu_result_13;
output 	W_alu_result_14;
output 	W_alu_result_15;
output 	W_alu_result_16;
output 	W_alu_result_3;
output 	W_alu_result_2;
output 	F_pc_9;
output 	F_pc_10;
output 	F_pc_11;
output 	F_pc_12;
output 	F_pc_14;
input 	q_a_22;
input 	q_a_23;
input 	q_a_11;
input 	q_a_12;
input 	q_a_13;
input 	q_a_14;
input 	q_a_15;
input 	q_a_16;
input 	q_a_1;
input 	q_a_3;
input 	q_a_4;
input 	q_a_5;
output 	F_pc_2;
input 	q_a_8;
input 	q_a_10;
input 	q_a_17;
output 	F_pc_8;
output 	F_pc_7;
output 	F_pc_6;
output 	F_pc_5;
output 	F_pc_4;
output 	F_pc_3;
input 	q_a_9;
input 	q_a_18;
input 	q_a_19;
input 	q_a_20;
input 	q_a_21;
output 	F_pc_1;
output 	F_pc_0;
output 	readdata_0;
output 	readdata_22;
output 	d_writedata_22;
output 	readdata_23;
output 	d_writedata_23;
output 	readdata_24;
output 	readdata_25;
output 	readdata_26;
output 	readdata_11;
output 	d_writedata_11;
output 	readdata_12;
output 	d_writedata_12;
output 	readdata_13;
output 	d_writedata_13;
output 	readdata_14;
output 	d_writedata_14;
output 	readdata_15;
output 	d_writedata_15;
output 	readdata_16;
output 	d_writedata_16;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_8;
output 	d_writedata_8;
output 	readdata_10;
output 	d_writedata_10;
output 	readdata_17;
output 	d_writedata_17;
output 	readdata_9;
output 	d_writedata_9;
output 	readdata_18;
output 	d_writedata_18;
output 	readdata_19;
output 	d_writedata_19;
output 	readdata_20;
output 	d_writedata_20;
output 	readdata_21;
output 	d_writedata_21;
input 	av_readdata_pre_16;
output 	readdata_6;
output 	readdata_7;
output 	readdata_27;
output 	readdata_28;
output 	readdata_29;
output 	readdata_30;
output 	readdata_31;
input 	av_readdata_pre_19;
input 	av_readdata_pre_18;
input 	av_readdata_pre_17;
input 	av_readdata_pre_20;
input 	av_readdata_pre_21;
input 	av_readdata_pre_22;
input 	av_waitrequest;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
output 	d_writedata_0;
input 	r_sync_rst;
output 	d_write1;
output 	d_writedata_1;
output 	d_writedata_2;
output 	d_writedata_3;
output 	d_writedata_4;
output 	d_writedata_5;
output 	d_read1;
input 	always2;
input 	av_waitrequest1;
input 	read_latency_shift_reg;
input 	saved_grant_0;
output 	debug_mem_slave_waitrequest;
input 	mem_used_1;
input 	WideOr0;
input 	src0_valid;
input 	read_latency_shift_reg_0;
input 	WideOr1;
input 	src1_valid;
output 	i_read1;
output 	F_pc_13;
input 	src_valid;
input 	mem;
output 	hbreak_enabled1;
input 	av_waitrequest2;
input 	src0_valid1;
input 	src_data_0;
input 	av_readdata_pre_221;
input 	src1_valid1;
input 	src1_valid2;
input 	src_data_22;
input 	av_readdata_pre_23;
input 	src_data_23;
input 	src_data_24;
input 	src_data_25;
input 	src_data_26;
input 	av_readdata_pre_11;
input 	av_readdata_pre_12;
input 	src_data_12;
input 	av_readdata_pre_13;
input 	av_readdata_pre_14;
input 	src_data_14;
input 	av_readdata_pre_15;
input 	av_readdata_pre_161;
input 	src_data_01;
input 	av_readdata_pre_1;
input 	src_data_2;
input 	av_readdata_pre_3;
input 	av_readdata_pre_4;
input 	av_readdata_pre_5;
input 	av_readdata_pre_8;
input 	src_data_8;
input 	av_readdata_pre_10;
input 	src_data_10;
input 	av_readdata_pre_171;
input 	src_data_17;
input 	av_readdata_pre_9;
input 	src_data_9;
input 	av_readdata_pre_181;
input 	av_readdata_pre_191;
input 	av_readdata_pre_201;
input 	av_readdata_pre_211;
input 	src_data_6;
input 	src_data_46;
input 	src_data_7;
input 	src_data_1;
input 	src_data_21;
input 	src_data_3;
input 	src_data_4;
input 	src_data_5;
input 	r_early_rst;
output 	d_byteenable_0;
input 	av_readdata_pre_81;
output 	d_byteenable_2;
output 	d_writedata_24;
output 	d_byteenable_3;
output 	d_writedata_25;
output 	d_writedata_26;
output 	d_byteenable_1;
input 	src_data_27;
input 	src_data_28;
input 	src_data_29;
input 	src_data_30;
input 	src_data_31;
input 	av_readdata_pre_101;
input 	av_readdata_pre_91;
input 	src_payload;
input 	src_payload1;
input 	av_readdata_pre_121;
input 	av_readdata_pre_131;
input 	av_readdata_pre_141;
input 	av_readdata_pre_151;
output 	d_writedata_6;
output 	d_writedata_7;
input 	src_payload2;
input 	src_data_38;
input 	src_data_41;
input 	src_data_45;
input 	src_data_44;
input 	src_data_43;
input 	src_data_42;
input 	src_data_40;
input 	src_data_39;
input 	src_payload3;
input 	src_data_32;
output 	d_writedata_27;
output 	d_writedata_28;
output 	d_writedata_29;
output 	d_writedata_30;
output 	d_writedata_31;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_data_34;
input 	src_payload16;
input 	src_payload17;
input 	src_data_35;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_data_33;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	src_payload33;
input 	src_payload34;
input 	src_payload35;
input 	src_payload36;
input 	src_payload37;
input 	src_payload38;
input 	src_payload39;
input 	src_payload40;
input 	src_payload41;
input 	src_payload42;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ;
wire \av_ld_byte0_data[0]~q ;
wire \W_alu_result[0]~q ;
wire \D_iw[22]~q ;
wire \D_iw[23]~q ;
wire \D_iw[24]~q ;
wire \D_iw[25]~q ;
wire \D_iw[26]~q ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ;
wire \av_ld_byte0_data[1]~q ;
wire \W_alu_result[1]~q ;
wire \av_ld_byte0_data[2]~q ;
wire \av_ld_byte0_data[3]~q ;
wire \av_ld_byte0_data[4]~q ;
wire \av_ld_byte0_data[5]~q ;
wire \W_estatus_reg~q ;
wire \D_iw[27]~q ;
wire \D_iw[28]~q ;
wire \D_iw[29]~q ;
wire \D_iw[30]~q ;
wire \D_iw[31]~q ;
wire \av_ld_byte0_data[7]~q ;
wire \av_ld_byte0_data[6]~q ;
wire \Add2~73_sumout ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ;
wire \niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ;
wire \av_ld_byte3_data[0]~q ;
wire \Add2~81_sumout ;
wire \av_ld_byte3_data[1]~q ;
wire \W_alu_result[25]~q ;
wire \av_ld_byte3_data[3]~q ;
wire \W_alu_result[27]~q ;
wire \W_alu_result[19]~q ;
wire \W_alu_result[20]~q ;
wire \W_alu_result[21]~q ;
wire \W_alu_result[22]~q ;
wire \W_alu_result[23]~q ;
wire \W_alu_result[24]~q ;
wire \W_alu_result[18]~q ;
wire \W_alu_result[17]~q ;
wire \av_ld_byte3_data[2]~q ;
wire \W_alu_result[26]~q ;
wire \av_ld_byte3_data[7]~q ;
wire \W_alu_result[31]~q ;
wire \av_ld_byte3_data[6]~q ;
wire \W_alu_result[30]~q ;
wire \av_ld_byte3_data[4]~q ;
wire \W_alu_result[28]~q ;
wire \av_ld_byte3_data[5]~q ;
wire \W_alu_result[29]~q ;
wire \Add2~85_sumout ;
wire \Add2~89_sumout ;
wire \Add2~93_sumout ;
wire \Add2~97_sumout ;
wire \Add2~101_sumout ;
wire \Add2~105_sumout ;
wire \Add2~109_sumout ;
wire \Add2~113_sumout ;
wire \Add2~117_sumout ;
wire \Add2~121_sumout ;
wire \Add2~125_sumout ;
wire \Add2~129_sumout ;
wire \Add2~133_sumout ;
wire \av_ld_byte2_data_nxt[6]~9_combout ;
wire \av_ld_byte2_data_nxt[5]~13_combout ;
wire \av_ld_byte2_data_nxt[4]~17_combout ;
wire \av_ld_byte2_data_nxt[1]~21_combout ;
wire \av_ld_byte2_data_nxt[2]~25_combout ;
wire \av_ld_byte2_data_nxt[3]~29_combout ;
wire \av_ld_byte2_data_nxt[0]~33_combout ;
wire \av_ld_byte1_data_nxt[7]~9_combout ;
wire \av_ld_byte1_data_nxt[6]~13_combout ;
wire \av_ld_byte1_data_nxt[5]~17_combout ;
wire \av_ld_byte1_data_nxt[4]~21_combout ;
wire \av_ld_byte1_data_nxt[1]~25_combout ;
wire \av_ld_byte1_data_nxt[2]~29_combout ;
wire \av_ld_byte1_data_nxt[0]~33_combout ;
wire \W_rf_wr_data[0]~31_combout ;
wire \R_wr_dst_reg~q ;
wire \W_rf_wren~combout ;
wire \W_control_rd_data[0]~q ;
wire \R_dst_regnum[0]~q ;
wire \R_dst_regnum[1]~q ;
wire \R_dst_regnum[2]~q ;
wire \R_dst_regnum[3]~q ;
wire \R_dst_regnum[4]~q ;
wire \W_rf_wr_data[1]~0_combout ;
wire \W_rf_wr_data[2]~1_combout ;
wire \W_rf_wr_data[3]~2_combout ;
wire \W_rf_wr_data[4]~3_combout ;
wire \W_rf_wr_data[5]~4_combout ;
wire \D_dst_regnum[1]~0_combout ;
wire \D_dst_regnum[1]~1_combout ;
wire \D_dst_regnum[2]~2_combout ;
wire \D_dst_regnum[2]~3_combout ;
wire \D_dst_regnum[0]~4_combout ;
wire \D_dst_regnum[0]~5_combout ;
wire \D_dst_regnum[3]~6_combout ;
wire \D_dst_regnum[3]~7_combout ;
wire \D_dst_regnum[4]~8_combout ;
wire \D_dst_regnum[4]~9_combout ;
wire \D_wr_dst_reg~0_combout ;
wire \D_wr_dst_reg~combout ;
wire \D_ctrl_ld_signed~0_combout ;
wire \av_ld_byte1_data[0]~q ;
wire \av_ld_rshift8~0_combout ;
wire \av_ld_byte0_data[2]~0_combout ;
wire \W_status_reg_pie~q ;
wire \Equal133~0_combout ;
wire \W_bstatus_reg~q ;
wire \E_control_rd_data[0]~0_combout ;
wire \E_alu_result[0]~16_combout ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci|the_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug|jtag_break~q ;
wire \av_ld_byte1_data[3]~q ;
wire \W_rf_wr_data[11]~5_combout ;
wire \av_ld_byte1_data[2]~q ;
wire \W_rf_wr_data[10]~6_combout ;
wire \av_ld_byte1_data[1]~q ;
wire \W_rf_wr_data[9]~7_combout ;
wire \W_rf_wr_data[8]~8_combout ;
wire \W_rf_wr_data[7]~9_combout ;
wire \W_rf_wr_data[6]~10_combout ;
wire \av_ld_byte1_data[4]~q ;
wire \W_rf_wr_data[12]~11_combout ;
wire \av_ld_byte1_data[5]~q ;
wire \W_rf_wr_data[13]~12_combout ;
wire \av_ld_byte1_data[6]~q ;
wire \W_rf_wr_data[14]~13_combout ;
wire \av_ld_byte1_data[7]~q ;
wire \W_rf_wr_data[15]~14_combout ;
wire \av_ld_byte2_data[0]~q ;
wire \W_rf_wr_data[16]~15_combout ;
wire \E_logic_result[1]~26_combout ;
wire \E_alu_result[1]~17_combout ;
wire \LessThan0~0_combout ;
wire \R_ctrl_ld_signed~q ;
wire \av_fill_bit~0_combout ;
wire \av_ld_byte1_data_en~0_combout ;
wire \R_ctrl_wrctl_inst~q ;
wire \W_status_reg_pie_inst_nxt~0_combout ;
wire \W_status_reg_pie_inst_nxt~1_combout ;
wire \W_status_reg_pie_inst_nxt~2_combout ;
wire \W_estatus_reg_inst_nxt~0_combout ;
wire \E_wrctl_bstatus~0_combout ;
wire \W_bstatus_reg_inst_nxt~0_combout ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci|the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_single_step_mode~q ;
wire \av_ld_byte2_data[3]~q ;
wire \av_ld_byte1_data_nxt[3]~0_combout ;
wire \av_ld_byte2_data[2]~q ;
wire \av_ld_byte2_data[1]~q ;
wire \av_ld_byte2_data[4]~q ;
wire \av_ld_byte2_data[5]~q ;
wire \av_ld_byte2_data[6]~q ;
wire \av_ld_byte2_data[7]~q ;
wire \W_rf_wr_data[25]~16_combout ;
wire \W_rf_wr_data[27]~17_combout ;
wire \W_rf_wr_data[19]~18_combout ;
wire \W_rf_wr_data[20]~19_combout ;
wire \W_rf_wr_data[21]~20_combout ;
wire \W_rf_wr_data[22]~21_combout ;
wire \W_rf_wr_data[23]~22_combout ;
wire \W_rf_wr_data[24]~23_combout ;
wire \W_rf_wr_data[18]~24_combout ;
wire \W_rf_wr_data[17]~25_combout ;
wire \W_rf_wr_data[26]~26_combout ;
wire \W_rf_wr_data[31]~27_combout ;
wire \W_rf_wr_data[30]~28_combout ;
wire \W_rf_wr_data[28]~29_combout ;
wire \W_rf_wr_data[29]~30_combout ;
wire \Equal62~17_combout ;
wire \D_op_wrctl~combout ;
wire \av_ld_byte2_data_nxt[7]~0_combout ;
wire \E_alu_result[25]~18_combout ;
wire \E_alu_result[27]~19_combout ;
wire \E_alu_result[19]~20_combout ;
wire \E_alu_result[20]~21_combout ;
wire \E_alu_result[21]~22_combout ;
wire \E_alu_result[22]~23_combout ;
wire \E_alu_result[23]~24_combout ;
wire \E_alu_result[24]~25_combout ;
wire \E_logic_result[18]~27_combout ;
wire \E_alu_result[18]~26_combout ;
wire \E_logic_result[17]~28_combout ;
wire \E_alu_result[17]~27_combout ;
wire \E_logic_result[26]~29_combout ;
wire \E_alu_result[26]~28_combout ;
wire \E_logic_result[31]~30_combout ;
wire \E_alu_result[31]~29_combout ;
wire \E_logic_result[30]~31_combout ;
wire \E_alu_result[30]~30_combout ;
wire \E_alu_result[28]~31_combout ;
wire \E_alu_result[29]~32_combout ;
wire \av_ld_byte1_data_nxt[3]~1_combout ;
wire \av_ld_byte2_data_nxt[7]~1_combout ;
wire \av_ld_byte1_data_nxt[0]~2_combout ;
wire \av_ld_byte1_data_nxt[2]~3_combout ;
wire \av_ld_byte1_data_nxt[1]~4_combout ;
wire \av_ld_byte1_data_nxt[4]~5_combout ;
wire \av_ld_byte1_data_nxt[5]~6_combout ;
wire \av_ld_byte1_data_nxt[6]~7_combout ;
wire \av_ld_byte1_data_nxt[7]~8_combout ;
wire \av_ld_byte2_data_nxt[0]~2_combout ;
wire \av_ld_byte2_data_nxt[3]~3_combout ;
wire \av_ld_byte2_data_nxt[2]~4_combout ;
wire \av_ld_byte2_data_nxt[1]~5_combout ;
wire \av_ld_byte2_data_nxt[4]~6_combout ;
wire \av_ld_byte2_data_nxt[5]~7_combout ;
wire \av_ld_byte2_data_nxt[6]~8_combout ;
wire \D_ctrl_implicit_dst_eretaddr~1_combout ;
wire \F_valid~0_combout ;
wire \D_valid~q ;
wire \R_valid~q ;
wire \E_new_inst~q ;
wire \D_iw[0]~q ;
wire \F_iw[1]~4_combout ;
wire \D_iw[1]~q ;
wire \F_iw[4]~6_combout ;
wire \D_iw[4]~q ;
wire \F_iw[3]~5_combout ;
wire \D_iw[3]~q ;
wire \D_ctrl_st~0_combout ;
wire \D_iw[2]~q ;
wire \R_ctrl_st~q ;
wire \d_write_nxt~0_combout ;
wire \D_ctrl_ld~0_combout ;
wire \R_ctrl_ld~q ;
wire \av_ld_waiting_for_data~q ;
wire \av_ld_waiting_for_data_nxt~0_combout ;
wire \D_ctrl_mem32~0_combout ;
wire \av_ld_aligning_data_nxt~1_combout ;
wire \av_ld_aligning_data_nxt~2_combout ;
wire \av_ld_aligning_data~q ;
wire \av_ld_align_cycle_nxt[0]~1_combout ;
wire \av_ld_align_cycle[0]~q ;
wire \av_ld_align_cycle_nxt[1]~0_combout ;
wire \av_ld_align_cycle[1]~q ;
wire \D_ctrl_mem16~0_combout ;
wire \av_ld_aligning_data_nxt~0_combout ;
wire \E_ld_stall~0_combout ;
wire \F_iw[5]~7_combout ;
wire \D_iw[5]~q ;
wire \D_ctrl_b_is_dst~0_combout ;
wire \R_ctrl_br_nxt~0_combout ;
wire \R_ctrl_br_nxt~1_combout ;
wire \R_ctrl_br_nxt~2_combout ;
wire \F_iw[13]~1_combout ;
wire \D_iw[13]~q ;
wire \D_iw[12]~q ;
wire \F_iw[15]~2_combout ;
wire \D_iw[15]~q ;
wire \F_iw[11]~0_combout ;
wire \D_iw[11]~q ;
wire \D_iw[14]~q ;
wire \Equal0~0_combout ;
wire \R_src2_use_imm~1_combout ;
wire \R_src2_use_imm~5_combout ;
wire \R_src2_use_imm~0_combout ;
wire \R_src2_use_imm~q ;
wire \D_ctrl_src_imm5_shift_rot~0_combout ;
wire \D_ctrl_src_imm5_shift_rot~1_combout ;
wire \R_ctrl_src_imm5_shift_rot~q ;
wire \R_src2_lo~0_combout ;
wire \D_ctrl_hi_imm16~0_combout ;
wire \R_ctrl_hi_imm16~q ;
wire \Equal62~7_combout ;
wire \Equal62~8_combout ;
wire \D_ctrl_implicit_dst_eretaddr~5_combout ;
wire \D_ctrl_implicit_dst_eretaddr~4_combout ;
wire \D_ctrl_implicit_dst_eretaddr~3_combout ;
wire \D_ctrl_implicit_dst_eretaddr~0_combout ;
wire \Equal0~10_combout ;
wire \D_ctrl_exception~6_combout ;
wire \D_ctrl_exception~5_combout ;
wire \D_ctrl_exception~4_combout ;
wire \D_ctrl_exception~1_combout ;
wire \Equal62~9_combout ;
wire \Equal62~10_combout ;
wire \Equal62~11_combout ;
wire \Equal62~13_combout ;
wire \Equal62~14_combout ;
wire \D_ctrl_force_src2_zero~0_combout ;
wire \Equal0~7_combout ;
wire \Equal0~8_combout ;
wire \D_ctrl_retaddr~2_combout ;
wire \D_ctrl_retaddr~0_combout ;
wire \Equal0~11_combout ;
wire \Equal62~15_combout ;
wire \Equal62~16_combout ;
wire \D_ctrl_force_src2_zero~1_combout ;
wire \D_ctrl_force_src2_zero~2_combout ;
wire \R_ctrl_force_src2_zero~q ;
wire \D_iw[6]~q ;
wire \R_src2_lo[0]~5_combout ;
wire \E_src2[0]~q ;
wire \E_shift_rot_cnt[0]~_wirecell_combout ;
wire \E_shift_rot_cnt[0]~q ;
wire \Add3~3_combout ;
wire \D_iw[7]~q ;
wire \R_src2_lo[1]~4_combout ;
wire \E_src2[1]~q ;
wire \E_shift_rot_cnt[1]~q ;
wire \Add3~2_combout ;
wire \D_iw[8]~q ;
wire \R_src2_lo[2]~3_combout ;
wire \E_src2[2]~q ;
wire \E_shift_rot_cnt[2]~q ;
wire \Add3~1_combout ;
wire \D_iw[9]~q ;
wire \R_src2_lo[3]~2_combout ;
wire \E_src2[3]~q ;
wire \E_shift_rot_cnt[3]~q ;
wire \E_shift_rot_done~0_combout ;
wire \Add3~0_combout ;
wire \D_iw[10]~q ;
wire \R_src2_lo[4]~1_combout ;
wire \E_src2[4]~q ;
wire \E_shift_rot_cnt[4]~q ;
wire \E_stall~0_combout ;
wire \E_stall~1_combout ;
wire \E_valid_from_R~0_combout ;
wire \E_valid_from_R~q ;
wire \W_valid~0_combout ;
wire \W_valid~q ;
wire \hbreak_pending_nxt~0_combout ;
wire \hbreak_pending~q ;
wire \wait_for_one_post_bret_inst~0_combout ;
wire \wait_for_one_post_bret_inst~q ;
wire \hbreak_req~0_combout ;
wire \F_iw[16]~3_combout ;
wire \D_iw[16]~q ;
wire \D_ctrl_shift_rot~0_combout ;
wire \D_ctrl_shift_rot~1_combout ;
wire \R_ctrl_shift_rot~q ;
wire \D_ctrl_shift_rot_right~0_combout ;
wire \D_ctrl_shift_rot_right~1_combout ;
wire \R_ctrl_shift_rot_right~q ;
wire \E_shift_rot_result_nxt[3]~13_combout ;
wire \R_ctrl_br~q ;
wire \D_ctrl_implicit_dst_eretaddr~2_combout ;
wire \Equal0~9_combout ;
wire \D_ctrl_retaddr~3_combout ;
wire \D_ctrl_retaddr~1_combout ;
wire \R_ctrl_retaddr~q ;
wire \R_src1~0_combout ;
wire \D_ctrl_jmp_direct~0_combout ;
wire \R_ctrl_jmp_direct~q ;
wire \R_src1~1_combout ;
wire \Add0~58 ;
wire \Add0~53_sumout ;
wire \R_src1[3]~15_combout ;
wire \E_src1[3]~q ;
wire \E_shift_rot_result[3]~q ;
wire \E_shift_rot_result_nxt[2]~14_combout ;
wire \Add0~57_sumout ;
wire \R_src1[2]~16_combout ;
wire \E_src1[2]~q ;
wire \E_shift_rot_result[2]~q ;
wire \E_shift_rot_result_nxt[1]~16_combout ;
wire \E_src1[26]~0_combout ;
wire \E_src1[1]~q ;
wire \E_shift_rot_result[1]~q ;
wire \E_shift_rot_result_nxt[0]~17_combout ;
wire \E_src1[0]~q ;
wire \E_shift_rot_result[0]~q ;
wire \Equal62~0_combout ;
wire \Equal62~2_combout ;
wire \D_ctrl_shift_logical~0_combout ;
wire \D_ctrl_shift_logical~1_combout ;
wire \R_ctrl_shift_logical~q ;
wire \Equal62~1_combout ;
wire \R_ctrl_rot_right_nxt~combout ;
wire \R_ctrl_rot_right~q ;
wire \E_shift_rot_fill_bit~0_combout ;
wire \E_shift_rot_result_nxt[31]~19_combout ;
wire \E_src1[31]~q ;
wire \E_shift_rot_result[31]~q ;
wire \E_shift_rot_result_nxt[30]~21_combout ;
wire \E_src1[30]~q ;
wire \E_shift_rot_result[30]~q ;
wire \E_shift_rot_result_nxt[29]~31_combout ;
wire \E_src1[29]~q ;
wire \E_shift_rot_result[29]~q ;
wire \E_shift_rot_result_nxt[28]~30_combout ;
wire \E_src1[28]~q ;
wire \E_shift_rot_result[28]~q ;
wire \E_shift_rot_result_nxt[27]~24_combout ;
wire \E_src1[27]~q ;
wire \E_shift_rot_result[27]~q ;
wire \E_shift_rot_result_nxt[26]~29_combout ;
wire \E_src1[26]~q ;
wire \E_shift_rot_result[26]~q ;
wire \E_shift_rot_result_nxt[25]~23_combout ;
wire \E_src1[25]~q ;
wire \E_shift_rot_result[25]~q ;
wire \E_shift_rot_result_nxt[24]~28_combout ;
wire \E_src1[24]~q ;
wire \E_shift_rot_result[24]~q ;
wire \E_shift_rot_result_nxt[23]~27_combout ;
wire \E_src1[23]~q ;
wire \E_shift_rot_result[23]~q ;
wire \E_shift_rot_result_nxt[22]~26_combout ;
wire \E_src1[22]~q ;
wire \E_shift_rot_result[22]~q ;
wire \E_shift_rot_result_nxt[21]~25_combout ;
wire \E_src1[21]~q ;
wire \E_shift_rot_result[21]~q ;
wire \E_shift_rot_result_nxt[20]~22_combout ;
wire \E_src1[20]~q ;
wire \E_shift_rot_result[20]~q ;
wire \E_shift_rot_result_nxt[19]~20_combout ;
wire \E_src1[19]~q ;
wire \E_shift_rot_result[19]~q ;
wire \E_shift_rot_result_nxt[18]~18_combout ;
wire \E_src1[18]~q ;
wire \E_shift_rot_result[18]~q ;
wire \E_shift_rot_result_nxt[17]~15_combout ;
wire \E_src1[17]~q ;
wire \E_shift_rot_result[17]~q ;
wire \E_shift_rot_result_nxt[16]~12_combout ;
wire \F_iw[20]~10_combout ;
wire \D_iw[20]~q ;
wire \Add0~54 ;
wire \Add0~2 ;
wire \Add0~30 ;
wire \Add0~26 ;
wire \Add0~22 ;
wire \Add0~18 ;
wire \Add0~14 ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~34 ;
wire \Add0~38 ;
wire \Add0~42 ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \R_src1[16]~14_combout ;
wire \E_src1[16]~q ;
wire \E_shift_rot_result[16]~q ;
wire \E_shift_rot_result_nxt[15]~11_combout ;
wire \F_iw[19]~9_combout ;
wire \D_iw[19]~q ;
wire \Add0~45_sumout ;
wire \R_src1[15]~13_combout ;
wire \E_src1[15]~q ;
wire \E_shift_rot_result[15]~q ;
wire \E_shift_rot_result_nxt[14]~10_combout ;
wire \F_iw[18]~8_combout ;
wire \D_iw[18]~q ;
wire \Add0~41_sumout ;
wire \R_src1[14]~12_combout ;
wire \E_src1[14]~q ;
wire \E_shift_rot_result[14]~q ;
wire \E_shift_rot_result_nxt[13]~9_combout ;
wire \D_iw[17]~q ;
wire \Add0~37_sumout ;
wire \R_src1[13]~11_combout ;
wire \E_src1[13]~q ;
wire \E_shift_rot_result[13]~q ;
wire \E_shift_rot_result_nxt[12]~8_combout ;
wire \Add0~33_sumout ;
wire \R_src1[12]~10_combout ;
wire \E_src1[12]~q ;
wire \E_shift_rot_result[12]~q ;
wire \E_shift_rot_result_nxt[11]~1_combout ;
wire \Add0~5_sumout ;
wire \R_src1[11]~3_combout ;
wire \E_src1[11]~q ;
wire \E_shift_rot_result[11]~q ;
wire \E_shift_rot_result_nxt[10]~2_combout ;
wire \Add0~9_sumout ;
wire \R_src1[10]~4_combout ;
wire \E_src1[10]~q ;
wire \E_shift_rot_result[10]~q ;
wire \E_shift_rot_result_nxt[9]~3_combout ;
wire \Add0~13_sumout ;
wire \R_src1[9]~5_combout ;
wire \E_src1[9]~q ;
wire \E_shift_rot_result[9]~q ;
wire \E_shift_rot_result_nxt[8]~4_combout ;
wire \Add0~17_sumout ;
wire \R_src1[8]~6_combout ;
wire \E_src1[8]~q ;
wire \E_shift_rot_result[8]~q ;
wire \E_shift_rot_result_nxt[7]~5_combout ;
wire \Add0~21_sumout ;
wire \R_src1[7]~7_combout ;
wire \E_src1[7]~q ;
wire \E_shift_rot_result[7]~q ;
wire \E_shift_rot_result_nxt[6]~6_combout ;
wire \Add0~25_sumout ;
wire \R_src1[6]~8_combout ;
wire \E_src1[6]~q ;
wire \E_shift_rot_result[6]~q ;
wire \E_shift_rot_result_nxt[5]~7_combout ;
wire \Add0~29_sumout ;
wire \R_src1[5]~9_combout ;
wire \E_src1[5]~q ;
wire \E_shift_rot_result[5]~q ;
wire \E_shift_rot_result_nxt[4]~0_combout ;
wire \Add0~1_sumout ;
wire \R_src1[4]~2_combout ;
wire \E_src1[4]~q ;
wire \E_shift_rot_result[4]~q ;
wire \D_ctrl_logic~0_combout ;
wire \D_ctrl_logic~1_combout ;
wire \R_ctrl_logic~q ;
wire \D_logic_op_raw[1]~0_combout ;
wire \D_ctrl_alu_force_xor~1_combout ;
wire \D_ctrl_alu_subtract~2_combout ;
wire \D_ctrl_alu_force_xor~0_combout ;
wire \D_logic_op[1]~0_combout ;
wire \R_logic_op[1]~q ;
wire \D_logic_op_raw[0]~1_combout ;
wire \D_logic_op[0]~1_combout ;
wire \R_logic_op[0]~q ;
wire \E_logic_result[4]~0_combout ;
wire \D_ctrl_alu_subtract~1_combout ;
wire \D_ctrl_alu_subtract~0_combout ;
wire \E_alu_sub~0_combout ;
wire \E_alu_sub~q ;
wire \Add2~78_cout ;
wire \Add2~70 ;
wire \Add2~62 ;
wire \Add2~58 ;
wire \Add2~54 ;
wire \Add2~1_sumout ;
wire \E_alu_result[4]~0_combout ;
wire \Equal62~4_combout ;
wire \D_op_rdctl~combout ;
wire \R_ctrl_rd_ctl_reg~q ;
wire \Equal62~5_combout ;
wire \Equal62~6_combout ;
wire \D_ctrl_unsigned_lo_imm16~1_combout ;
wire \Equal0~1_combout ;
wire \Equal0~4_combout ;
wire \Equal0~5_combout ;
wire \Equal0~6_combout ;
wire \D_ctrl_br_cmp~0_combout ;
wire \D_ctrl_br_cmp~1_combout ;
wire \R_ctrl_br_cmp~q ;
wire \E_alu_result~1_combout ;
wire \E_src2[15]~0_combout ;
wire \E_src2[11]~q ;
wire \E_logic_result[11]~1_combout ;
wire \E_src2[10]~q ;
wire \E_src2[9]~q ;
wire \E_src2[8]~q ;
wire \E_src2[7]~q ;
wire \E_src2[6]~q ;
wire \E_src2[5]~q ;
wire \Add2~2 ;
wire \Add2~30 ;
wire \Add2~26 ;
wire \Add2~22 ;
wire \Add2~18 ;
wire \Add2~14 ;
wire \Add2~10 ;
wire \Add2~5_sumout ;
wire \E_alu_result[11]~2_combout ;
wire \E_logic_result[10]~2_combout ;
wire \Add2~9_sumout ;
wire \E_alu_result[10]~3_combout ;
wire \E_logic_result[9]~3_combout ;
wire \Add2~13_sumout ;
wire \E_alu_result[9]~4_combout ;
wire \E_logic_result[8]~4_combout ;
wire \Add2~17_sumout ;
wire \E_alu_result[8]~5_combout ;
wire \E_logic_result[7]~5_combout ;
wire \Add2~21_sumout ;
wire \E_alu_result[7]~6_combout ;
wire \E_logic_result[6]~6_combout ;
wire \Add2~25_sumout ;
wire \E_alu_result[6]~7_combout ;
wire \E_logic_result[5]~7_combout ;
wire \Add2~29_sumout ;
wire \E_alu_result[5]~8_combout ;
wire \E_src2[12]~q ;
wire \E_logic_result[12]~8_combout ;
wire \Add2~6 ;
wire \Add2~33_sumout ;
wire \E_alu_result[12]~9_combout ;
wire \E_src2[13]~q ;
wire \E_logic_result[13]~9_combout ;
wire \Add2~34 ;
wire \Add2~37_sumout ;
wire \E_alu_result[13]~10_combout ;
wire \E_src2[14]~q ;
wire \E_logic_result[14]~10_combout ;
wire \Add2~38 ;
wire \Add2~41_sumout ;
wire \E_alu_result[14]~11_combout ;
wire \F_iw[21]~11_combout ;
wire \D_iw[21]~q ;
wire \E_src2[15]~q ;
wire \E_logic_result[15]~11_combout ;
wire \Add2~42 ;
wire \Add2~45_sumout ;
wire \E_alu_result[15]~12_combout ;
wire \R_src2_hi[0]~0_combout ;
wire \D_ctrl_logic~2_combout ;
wire \D_ctrl_unsigned_lo_imm16~0_combout ;
wire \R_ctrl_unsigned_lo_imm16~q ;
wire \R_src2_hi~1_combout ;
wire \E_src2[16]~q ;
wire \E_logic_result[16]~12_combout ;
wire \Add2~46 ;
wire \Add2~49_sumout ;
wire \E_alu_result[16]~13_combout ;
wire \E_logic_result[3]~13_combout ;
wire \Add2~53_sumout ;
wire \E_alu_result[3]~14_combout ;
wire \E_logic_result[2]~14_combout ;
wire \Add2~57_sumout ;
wire \E_alu_result[2]~15_combout ;
wire \D_ctrl_exception~0_combout ;
wire \D_ctrl_exception~3_combout ;
wire \D_ctrl_exception~2_combout ;
wire \R_ctrl_exception~q ;
wire \D_ctrl_break~0_combout ;
wire \R_ctrl_break~q ;
wire \F_pc_sel_nxt.01~0_combout ;
wire \Equal0~12_combout ;
wire \Equal62~3_combout ;
wire \Equal0~2_combout ;
wire \E_invert_arith_src_msb~0_combout ;
wire \E_invert_arith_src_msb~1_combout ;
wire \E_invert_arith_src_msb~q ;
wire \R_src2_hi[15]~13_combout ;
wire \E_src2[31]~q ;
wire \R_src2_hi[14]~14_combout ;
wire \E_src2[30]~q ;
wire \R_src2_hi[13]~16_combout ;
wire \E_src2[29]~q ;
wire \R_src2_hi[12]~15_combout ;
wire \E_src2[28]~q ;
wire \R_src2_hi[11]~3_combout ;
wire \E_src2[27]~q ;
wire \R_src2_hi[10]~12_combout ;
wire \E_src2[26]~q ;
wire \R_src2_hi[9]~2_combout ;
wire \E_src2[25]~q ;
wire \R_src2_hi[8]~9_combout ;
wire \E_src2[24]~q ;
wire \R_src2_hi[7]~8_combout ;
wire \E_src2[23]~q ;
wire \R_src2_hi[6]~7_combout ;
wire \E_src2[22]~q ;
wire \R_src2_hi[5]~6_combout ;
wire \E_src2[21]~q ;
wire \R_src2_hi[4]~5_combout ;
wire \E_src2[20]~q ;
wire \R_src2_hi[3]~4_combout ;
wire \E_src2[19]~q ;
wire \R_src2_hi[2]~10_combout ;
wire \E_src2[18]~q ;
wire \R_src2_hi[1]~11_combout ;
wire \E_src2[17]~q ;
wire \Add2~50 ;
wire \Add2~126 ;
wire \Add2~122 ;
wire \Add2~98 ;
wire \Add2~102 ;
wire \Add2~106 ;
wire \Add2~110 ;
wire \Add2~114 ;
wire \Add2~118 ;
wire \Add2~90 ;
wire \Add2~130 ;
wire \Add2~94 ;
wire \Add2~134 ;
wire \Add2~86 ;
wire \Add2~82 ;
wire \Add2~74 ;
wire \Add2~65_sumout ;
wire \R_compare_op[0]~q ;
wire \E_logic_result[25]~15_combout ;
wire \E_logic_result[27]~16_combout ;
wire \Equal127~0_combout ;
wire \E_logic_result[19]~17_combout ;
wire \E_logic_result[20]~18_combout ;
wire \E_logic_result[21]~19_combout ;
wire \E_logic_result[22]~20_combout ;
wire \E_logic_result[23]~21_combout ;
wire \E_logic_result[24]~22_combout ;
wire \Equal127~1_combout ;
wire \Equal127~2_combout ;
wire \Equal127~3_combout ;
wire \Equal127~4_combout ;
wire \Equal127~5_combout ;
wire \Equal127~6_combout ;
wire \Equal127~7_combout ;
wire \Equal127~8_combout ;
wire \Equal127~9_combout ;
wire \Equal127~10_combout ;
wire \E_logic_result[0]~23_combout ;
wire \E_logic_result[28]~24_combout ;
wire \E_logic_result[29]~25_combout ;
wire \Equal127~11_combout ;
wire \Equal127~12_combout ;
wire \R_compare_op[1]~q ;
wire \E_cmp_result~0_combout ;
wire \W_cmp_result~q ;
wire \Equal62~12_combout ;
wire \D_ctrl_uncond_cti_non_br~0_combout ;
wire \D_ctrl_uncond_cti_non_br~1_combout ;
wire \R_ctrl_uncond_cti_non_br~q ;
wire \Equal0~3_combout ;
wire \R_ctrl_br_uncond~q ;
wire \F_pc_sel_nxt~0_combout ;
wire \F_pc_sel_nxt.10~0_combout ;
wire \F_pc_no_crst_nxt[9]~0_combout ;
wire \F_pc_no_crst_nxt[10]~1_combout ;
wire \F_pc_no_crst_nxt[11]~2_combout ;
wire \F_pc_no_crst_nxt[12]~3_combout ;
wire \F_pc_no_crst_nxt[14]~5_combout ;
wire \F_pc_no_crst_nxt[2]~6_combout ;
wire \F_pc_no_crst_nxt[8]~7_combout ;
wire \F_pc_no_crst_nxt[7]~8_combout ;
wire \F_pc_no_crst_nxt[6]~9_combout ;
wire \F_pc_no_crst_nxt[5]~10_combout ;
wire \F_pc_no_crst_nxt[4]~11_combout ;
wire \F_pc_no_crst_nxt~12_combout ;
wire \F_pc_no_crst_nxt[1]~13_combout ;
wire \F_pc_no_crst_nxt[0]~14_combout ;
wire \D_ctrl_mem8~0_combout ;
wire \E_st_data[23]~0_combout ;
wire \D_ctrl_mem8~1_combout ;
wire \E_st_stall~combout ;
wire \d_read_nxt~combout ;
wire \i_read_nxt~0_combout ;
wire \F_pc_no_crst_nxt[13]~4_combout ;
wire \hbreak_enabled~0_combout ;
wire \Add2~61_sumout ;
wire \D_ctrl_mem16~1_combout ;
wire \Add2~69_sumout ;
wire \E_mem_byte_en~0_combout ;
wire \E_mem_byte_en[2]~1_combout ;
wire \E_st_data[24]~1_combout ;
wire \E_mem_byte_en[3]~2_combout ;
wire \E_st_data[25]~2_combout ;
wire \E_st_data[26]~3_combout ;
wire \E_mem_byte_en[1]~3_combout ;
wire \E_st_data[27]~4_combout ;
wire \E_st_data[28]~5_combout ;
wire \E_st_data[29]~6_combout ;
wire \E_st_data[30]~7_combout ;
wire \E_st_data[31]~8_combout ;


niosLab2_niosLab2_nios2_gen2_0_cpu_register_bank_b_module niosLab2_nios2_gen2_0_cpu_register_bank_b(
	.q_b_0(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_1(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_2(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_3(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_4(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_5(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.D_iw_22(\D_iw[22]~q ),
	.D_iw_23(\D_iw[23]~q ),
	.D_iw_24(\D_iw[24]~q ),
	.D_iw_25(\D_iw[25]~q ),
	.D_iw_26(\D_iw[26]~q ),
	.q_b_11(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_7(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_6(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_12(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_13(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_14(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_15(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_16(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_25(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_27(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_19(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_20(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_21(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_22(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_23(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_24(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_18(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_17(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_26(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_31(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_30(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_28(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_29(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.W_rf_wr_data_0(\W_rf_wr_data[0]~31_combout ),
	.W_rf_wren(\W_rf_wren~combout ),
	.R_dst_regnum_0(\R_dst_regnum[0]~q ),
	.R_dst_regnum_1(\R_dst_regnum[1]~q ),
	.R_dst_regnum_2(\R_dst_regnum[2]~q ),
	.R_dst_regnum_3(\R_dst_regnum[3]~q ),
	.R_dst_regnum_4(\R_dst_regnum[4]~q ),
	.W_rf_wr_data_1(\W_rf_wr_data[1]~0_combout ),
	.W_rf_wr_data_2(\W_rf_wr_data[2]~1_combout ),
	.W_rf_wr_data_3(\W_rf_wr_data[3]~2_combout ),
	.W_rf_wr_data_4(\W_rf_wr_data[4]~3_combout ),
	.W_rf_wr_data_5(\W_rf_wr_data[5]~4_combout ),
	.W_rf_wr_data_11(\W_rf_wr_data[11]~5_combout ),
	.W_rf_wr_data_10(\W_rf_wr_data[10]~6_combout ),
	.W_rf_wr_data_9(\W_rf_wr_data[9]~7_combout ),
	.W_rf_wr_data_8(\W_rf_wr_data[8]~8_combout ),
	.W_rf_wr_data_7(\W_rf_wr_data[7]~9_combout ),
	.W_rf_wr_data_6(\W_rf_wr_data[6]~10_combout ),
	.W_rf_wr_data_12(\W_rf_wr_data[12]~11_combout ),
	.W_rf_wr_data_13(\W_rf_wr_data[13]~12_combout ),
	.W_rf_wr_data_14(\W_rf_wr_data[14]~13_combout ),
	.W_rf_wr_data_15(\W_rf_wr_data[15]~14_combout ),
	.W_rf_wr_data_16(\W_rf_wr_data[16]~15_combout ),
	.W_rf_wr_data_25(\W_rf_wr_data[25]~16_combout ),
	.W_rf_wr_data_27(\W_rf_wr_data[27]~17_combout ),
	.W_rf_wr_data_19(\W_rf_wr_data[19]~18_combout ),
	.W_rf_wr_data_20(\W_rf_wr_data[20]~19_combout ),
	.W_rf_wr_data_21(\W_rf_wr_data[21]~20_combout ),
	.W_rf_wr_data_22(\W_rf_wr_data[22]~21_combout ),
	.W_rf_wr_data_23(\W_rf_wr_data[23]~22_combout ),
	.W_rf_wr_data_24(\W_rf_wr_data[24]~23_combout ),
	.W_rf_wr_data_18(\W_rf_wr_data[18]~24_combout ),
	.W_rf_wr_data_17(\W_rf_wr_data[17]~25_combout ),
	.W_rf_wr_data_26(\W_rf_wr_data[26]~26_combout ),
	.W_rf_wr_data_31(\W_rf_wr_data[31]~27_combout ),
	.W_rf_wr_data_30(\W_rf_wr_data[30]~28_combout ),
	.W_rf_wr_data_28(\W_rf_wr_data[28]~29_combout ),
	.W_rf_wr_data_29(\W_rf_wr_data[29]~30_combout ),
	.clk_clk(clk_clk));

niosLab2_niosLab2_nios2_gen2_0_cpu_register_bank_a_module niosLab2_nios2_gen2_0_cpu_register_bank_a(
	.q_b_4(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_11(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_7(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_6(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_5(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_12(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_13(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_14(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_15(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_16(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_3(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_2(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.D_iw_27(\D_iw[27]~q ),
	.D_iw_28(\D_iw[28]~q ),
	.D_iw_29(\D_iw[29]~q ),
	.D_iw_30(\D_iw[30]~q ),
	.D_iw_31(\D_iw[31]~q ),
	.q_b_25(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_27(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_19(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_20(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_21(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_22(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_23(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_24(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_18(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_17(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_1(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_26(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_31(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_30(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_0(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_28(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_29(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.W_rf_wr_data_0(\W_rf_wr_data[0]~31_combout ),
	.W_rf_wren(\W_rf_wren~combout ),
	.R_dst_regnum_0(\R_dst_regnum[0]~q ),
	.R_dst_regnum_1(\R_dst_regnum[1]~q ),
	.R_dst_regnum_2(\R_dst_regnum[2]~q ),
	.R_dst_regnum_3(\R_dst_regnum[3]~q ),
	.R_dst_regnum_4(\R_dst_regnum[4]~q ),
	.W_rf_wr_data_1(\W_rf_wr_data[1]~0_combout ),
	.W_rf_wr_data_2(\W_rf_wr_data[2]~1_combout ),
	.W_rf_wr_data_3(\W_rf_wr_data[3]~2_combout ),
	.W_rf_wr_data_4(\W_rf_wr_data[4]~3_combout ),
	.W_rf_wr_data_5(\W_rf_wr_data[5]~4_combout ),
	.W_rf_wr_data_11(\W_rf_wr_data[11]~5_combout ),
	.W_rf_wr_data_10(\W_rf_wr_data[10]~6_combout ),
	.W_rf_wr_data_9(\W_rf_wr_data[9]~7_combout ),
	.W_rf_wr_data_8(\W_rf_wr_data[8]~8_combout ),
	.W_rf_wr_data_7(\W_rf_wr_data[7]~9_combout ),
	.W_rf_wr_data_6(\W_rf_wr_data[6]~10_combout ),
	.W_rf_wr_data_12(\W_rf_wr_data[12]~11_combout ),
	.W_rf_wr_data_13(\W_rf_wr_data[13]~12_combout ),
	.W_rf_wr_data_14(\W_rf_wr_data[14]~13_combout ),
	.W_rf_wr_data_15(\W_rf_wr_data[15]~14_combout ),
	.W_rf_wr_data_16(\W_rf_wr_data[16]~15_combout ),
	.W_rf_wr_data_25(\W_rf_wr_data[25]~16_combout ),
	.W_rf_wr_data_27(\W_rf_wr_data[27]~17_combout ),
	.W_rf_wr_data_19(\W_rf_wr_data[19]~18_combout ),
	.W_rf_wr_data_20(\W_rf_wr_data[20]~19_combout ),
	.W_rf_wr_data_21(\W_rf_wr_data[21]~20_combout ),
	.W_rf_wr_data_22(\W_rf_wr_data[22]~21_combout ),
	.W_rf_wr_data_23(\W_rf_wr_data[23]~22_combout ),
	.W_rf_wr_data_24(\W_rf_wr_data[24]~23_combout ),
	.W_rf_wr_data_18(\W_rf_wr_data[18]~24_combout ),
	.W_rf_wr_data_17(\W_rf_wr_data[17]~25_combout ),
	.W_rf_wr_data_26(\W_rf_wr_data[26]~26_combout ),
	.W_rf_wr_data_31(\W_rf_wr_data[31]~27_combout ),
	.W_rf_wr_data_30(\W_rf_wr_data[30]~28_combout ),
	.W_rf_wr_data_28(\W_rf_wr_data[28]~29_combout ),
	.W_rf_wr_data_29(\W_rf_wr_data[29]~30_combout ),
	.clk_clk(clk_clk));

niosLab2_niosLab2_nios2_gen2_0_cpu_nios2_oci the_niosLab2_nios2_gen2_0_cpu_nios2_oci(
	.readdata_0(readdata_0),
	.readdata_22(readdata_22),
	.readdata_23(readdata_23),
	.readdata_24(readdata_24),
	.readdata_25(readdata_25),
	.readdata_26(readdata_26),
	.readdata_11(readdata_11),
	.readdata_12(readdata_12),
	.readdata_13(readdata_13),
	.readdata_14(readdata_14),
	.readdata_15(readdata_15),
	.readdata_16(readdata_16),
	.readdata_1(readdata_1),
	.readdata_2(readdata_2),
	.readdata_3(readdata_3),
	.readdata_4(readdata_4),
	.readdata_5(readdata_5),
	.readdata_8(readdata_8),
	.readdata_10(readdata_10),
	.readdata_17(readdata_17),
	.readdata_9(readdata_9),
	.readdata_18(readdata_18),
	.readdata_19(readdata_19),
	.readdata_20(readdata_20),
	.readdata_21(readdata_21),
	.readdata_6(readdata_6),
	.readdata_7(readdata_7),
	.readdata_27(readdata_27),
	.readdata_28(readdata_28),
	.readdata_29(readdata_29),
	.readdata_30(readdata_30),
	.readdata_31(readdata_31),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.r_sync_rst(r_sync_rst),
	.always2(always2),
	.saved_grant_0(saved_grant_0),
	.waitrequest(debug_mem_slave_waitrequest),
	.mem_used_1(mem_used_1),
	.src1_valid(src1_valid),
	.src_valid(src_valid),
	.mem(mem),
	.hbreak_enabled(hbreak_enabled1),
	.jtag_break(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci|the_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug|jtag_break~q ),
	.address_nxt({src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.r_early_rst(r_early_rst),
	.oci_single_step_mode(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci|the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.writedata_nxt({src_payload42,src_payload41,src_payload40,src_payload39,src_payload38,src_payload19,src_payload18,src_payload17,src_payload16,src_payload15,src_payload35,src_payload34,src_payload33,src_payload32,src_payload30,src_payload25,src_payload24,src_payload23,src_payload22,
src_payload21,src_payload20,src_payload29,src_payload31,src_payload28,src_payload37,src_payload36,src_payload27,src_payload26,src_payload13,src_payload14,src_payload5,src_payload2}),
	.debugaccess_nxt(src_payload3),
	.byteenable_nxt({src_data_35,src_data_34,src_data_33,src_data_32}),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

dffeas \av_ld_byte0_data[0] (
	.clk(clk_clk),
	.d(src_data_0),
	.asdata(\av_ld_byte1_data[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~0_combout ),
	.ena(\av_ld_byte0_data[2]~0_combout ),
	.q(\av_ld_byte0_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[0] .power_up = "low";

dffeas \W_alu_result[0] (
	.clk(clk_clk),
	.d(\E_alu_result[0]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[0]~q ),
	.prn(vcc));
defparam \W_alu_result[0] .is_wysiwyg = "true";
defparam \W_alu_result[0] .power_up = "low";

dffeas \D_iw[22] (
	.clk(clk_clk),
	.d(src_data_22),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[22]~q ),
	.prn(vcc));
defparam \D_iw[22] .is_wysiwyg = "true";
defparam \D_iw[22] .power_up = "low";

dffeas \D_iw[23] (
	.clk(clk_clk),
	.d(src_data_23),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[23]~q ),
	.prn(vcc));
defparam \D_iw[23] .is_wysiwyg = "true";
defparam \D_iw[23] .power_up = "low";

dffeas \D_iw[24] (
	.clk(clk_clk),
	.d(src_data_24),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[24]~q ),
	.prn(vcc));
defparam \D_iw[24] .is_wysiwyg = "true";
defparam \D_iw[24] .power_up = "low";

dffeas \D_iw[25] (
	.clk(clk_clk),
	.d(src_data_25),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[25]~q ),
	.prn(vcc));
defparam \D_iw[25] .is_wysiwyg = "true";
defparam \D_iw[25] .power_up = "low";

dffeas \D_iw[26] (
	.clk(clk_clk),
	.d(src_data_26),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[26]~q ),
	.prn(vcc));
defparam \D_iw[26] .is_wysiwyg = "true";
defparam \D_iw[26] .power_up = "low";

dffeas \av_ld_byte0_data[1] (
	.clk(clk_clk),
	.d(src_data_1),
	.asdata(\av_ld_byte1_data[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~0_combout ),
	.ena(\av_ld_byte0_data[2]~0_combout ),
	.q(\av_ld_byte0_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[1] .power_up = "low";

dffeas \W_alu_result[1] (
	.clk(clk_clk),
	.d(\E_alu_result[1]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[1]~q ),
	.prn(vcc));
defparam \W_alu_result[1] .is_wysiwyg = "true";
defparam \W_alu_result[1] .power_up = "low";

dffeas \av_ld_byte0_data[2] (
	.clk(clk_clk),
	.d(src_data_21),
	.asdata(\av_ld_byte1_data[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~0_combout ),
	.ena(\av_ld_byte0_data[2]~0_combout ),
	.q(\av_ld_byte0_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[2] .power_up = "low";

dffeas \av_ld_byte0_data[3] (
	.clk(clk_clk),
	.d(src_data_3),
	.asdata(\av_ld_byte1_data[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~0_combout ),
	.ena(\av_ld_byte0_data[2]~0_combout ),
	.q(\av_ld_byte0_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[3] .power_up = "low";

dffeas \av_ld_byte0_data[4] (
	.clk(clk_clk),
	.d(src_data_4),
	.asdata(\av_ld_byte1_data[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~0_combout ),
	.ena(\av_ld_byte0_data[2]~0_combout ),
	.q(\av_ld_byte0_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[4] .power_up = "low";

dffeas \av_ld_byte0_data[5] (
	.clk(clk_clk),
	.d(src_data_5),
	.asdata(\av_ld_byte1_data[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~0_combout ),
	.ena(\av_ld_byte0_data[2]~0_combout ),
	.q(\av_ld_byte0_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[5] .power_up = "low";

dffeas W_estatus_reg(
	.clk(clk_clk),
	.d(\W_estatus_reg_inst_nxt~0_combout ),
	.asdata(\W_status_reg_pie~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_ctrl_exception~q ),
	.ena(\E_valid_from_R~q ),
	.q(\W_estatus_reg~q ),
	.prn(vcc));
defparam W_estatus_reg.is_wysiwyg = "true";
defparam W_estatus_reg.power_up = "low";

dffeas \D_iw[27] (
	.clk(clk_clk),
	.d(src_data_27),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[27]~q ),
	.prn(vcc));
defparam \D_iw[27] .is_wysiwyg = "true";
defparam \D_iw[27] .power_up = "low";

dffeas \D_iw[28] (
	.clk(clk_clk),
	.d(src_data_28),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[28]~q ),
	.prn(vcc));
defparam \D_iw[28] .is_wysiwyg = "true";
defparam \D_iw[28] .power_up = "low";

dffeas \D_iw[29] (
	.clk(clk_clk),
	.d(src_data_29),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[29]~q ),
	.prn(vcc));
defparam \D_iw[29] .is_wysiwyg = "true";
defparam \D_iw[29] .power_up = "low";

dffeas \D_iw[30] (
	.clk(clk_clk),
	.d(src_data_30),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[30]~q ),
	.prn(vcc));
defparam \D_iw[30] .is_wysiwyg = "true";
defparam \D_iw[30] .power_up = "low";

dffeas \D_iw[31] (
	.clk(clk_clk),
	.d(src_data_31),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[31]~q ),
	.prn(vcc));
defparam \D_iw[31] .is_wysiwyg = "true";
defparam \D_iw[31] .power_up = "low";

dffeas \av_ld_byte0_data[7] (
	.clk(clk_clk),
	.d(src_payload),
	.asdata(\av_ld_byte1_data[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~0_combout ),
	.ena(\av_ld_byte0_data[2]~0_combout ),
	.q(\av_ld_byte0_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[7] .power_up = "low";

dffeas \av_ld_byte0_data[6] (
	.clk(clk_clk),
	.d(src_payload1),
	.asdata(\av_ld_byte1_data[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~0_combout ),
	.ena(\av_ld_byte0_data[2]~0_combout ),
	.q(\av_ld_byte0_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[6] .power_up = "low";

cyclonev_lcell_comb \Add2~73 (
	.dataa(!\E_invert_arith_src_msb~q ),
	.datab(!\E_alu_sub~q ),
	.datac(gnd),
	.datad(!\E_src2[31]~q ),
	.datae(gnd),
	.dataf(!\E_src1[31]~q ),
	.datag(gnd),
	.cin(\Add2~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~73_sumout ),
	.cout(\Add2~74 ),
	.shareout());
defparam \Add2~73 .extended_lut = "off";
defparam \Add2~73 .lut_mask = 64'h000055AA00009966;
defparam \Add2~73 .shared_arith = "off";

dffeas \av_ld_byte3_data[0] (
	.clk(clk_clk),
	.d(src_payload4),
	.asdata(\av_fill_bit~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_aligning_data~q ),
	.ena(!\av_ld_rshift8~0_combout ),
	.q(\av_ld_byte3_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[0] .power_up = "low";

cyclonev_lcell_comb \Add2~81 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[30]~q ),
	.datae(gnd),
	.dataf(!\E_src1[30]~q ),
	.datag(gnd),
	.cin(\Add2~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~81_sumout ),
	.cout(\Add2~82 ),
	.shareout());
defparam \Add2~81 .extended_lut = "off";
defparam \Add2~81 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~81 .shared_arith = "off";

dffeas \av_ld_byte3_data[1] (
	.clk(clk_clk),
	.d(src_payload6),
	.asdata(\av_fill_bit~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_aligning_data~q ),
	.ena(!\av_ld_rshift8~0_combout ),
	.q(\av_ld_byte3_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[1] .power_up = "low";

dffeas \W_alu_result[25] (
	.clk(clk_clk),
	.d(\E_alu_result[25]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[25]~q ),
	.prn(vcc));
defparam \W_alu_result[25] .is_wysiwyg = "true";
defparam \W_alu_result[25] .power_up = "low";

dffeas \av_ld_byte3_data[3] (
	.clk(clk_clk),
	.d(src_payload7),
	.asdata(\av_fill_bit~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_aligning_data~q ),
	.ena(!\av_ld_rshift8~0_combout ),
	.q(\av_ld_byte3_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[3] .power_up = "low";

dffeas \W_alu_result[27] (
	.clk(clk_clk),
	.d(\E_alu_result[27]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[27]~q ),
	.prn(vcc));
defparam \W_alu_result[27] .is_wysiwyg = "true";
defparam \W_alu_result[27] .power_up = "low";

dffeas \W_alu_result[19] (
	.clk(clk_clk),
	.d(\E_alu_result[19]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[19]~q ),
	.prn(vcc));
defparam \W_alu_result[19] .is_wysiwyg = "true";
defparam \W_alu_result[19] .power_up = "low";

dffeas \W_alu_result[20] (
	.clk(clk_clk),
	.d(\E_alu_result[20]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[20]~q ),
	.prn(vcc));
defparam \W_alu_result[20] .is_wysiwyg = "true";
defparam \W_alu_result[20] .power_up = "low";

dffeas \W_alu_result[21] (
	.clk(clk_clk),
	.d(\E_alu_result[21]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[21]~q ),
	.prn(vcc));
defparam \W_alu_result[21] .is_wysiwyg = "true";
defparam \W_alu_result[21] .power_up = "low";

dffeas \W_alu_result[22] (
	.clk(clk_clk),
	.d(\E_alu_result[22]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[22]~q ),
	.prn(vcc));
defparam \W_alu_result[22] .is_wysiwyg = "true";
defparam \W_alu_result[22] .power_up = "low";

dffeas \W_alu_result[23] (
	.clk(clk_clk),
	.d(\E_alu_result[23]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[23]~q ),
	.prn(vcc));
defparam \W_alu_result[23] .is_wysiwyg = "true";
defparam \W_alu_result[23] .power_up = "low";

dffeas \W_alu_result[24] (
	.clk(clk_clk),
	.d(\E_alu_result[24]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[24]~q ),
	.prn(vcc));
defparam \W_alu_result[24] .is_wysiwyg = "true";
defparam \W_alu_result[24] .power_up = "low";

dffeas \W_alu_result[18] (
	.clk(clk_clk),
	.d(\E_alu_result[18]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[18]~q ),
	.prn(vcc));
defparam \W_alu_result[18] .is_wysiwyg = "true";
defparam \W_alu_result[18] .power_up = "low";

dffeas \W_alu_result[17] (
	.clk(clk_clk),
	.d(\E_alu_result[17]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[17]~q ),
	.prn(vcc));
defparam \W_alu_result[17] .is_wysiwyg = "true";
defparam \W_alu_result[17] .power_up = "low";

dffeas \av_ld_byte3_data[2] (
	.clk(clk_clk),
	.d(src_payload8),
	.asdata(\av_fill_bit~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_aligning_data~q ),
	.ena(!\av_ld_rshift8~0_combout ),
	.q(\av_ld_byte3_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[2] .power_up = "low";

dffeas \W_alu_result[26] (
	.clk(clk_clk),
	.d(\E_alu_result[26]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[26]~q ),
	.prn(vcc));
defparam \W_alu_result[26] .is_wysiwyg = "true";
defparam \W_alu_result[26] .power_up = "low";

dffeas \av_ld_byte3_data[7] (
	.clk(clk_clk),
	.d(src_payload9),
	.asdata(\av_fill_bit~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_aligning_data~q ),
	.ena(!\av_ld_rshift8~0_combout ),
	.q(\av_ld_byte3_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[7] .power_up = "low";

dffeas \W_alu_result[31] (
	.clk(clk_clk),
	.d(\E_alu_result[31]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[31]~q ),
	.prn(vcc));
defparam \W_alu_result[31] .is_wysiwyg = "true";
defparam \W_alu_result[31] .power_up = "low";

dffeas \av_ld_byte3_data[6] (
	.clk(clk_clk),
	.d(src_payload10),
	.asdata(\av_fill_bit~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_aligning_data~q ),
	.ena(!\av_ld_rshift8~0_combout ),
	.q(\av_ld_byte3_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[6] .power_up = "low";

dffeas \W_alu_result[30] (
	.clk(clk_clk),
	.d(\E_alu_result[30]~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[30]~q ),
	.prn(vcc));
defparam \W_alu_result[30] .is_wysiwyg = "true";
defparam \W_alu_result[30] .power_up = "low";

dffeas \av_ld_byte3_data[4] (
	.clk(clk_clk),
	.d(src_payload11),
	.asdata(\av_fill_bit~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_aligning_data~q ),
	.ena(!\av_ld_rshift8~0_combout ),
	.q(\av_ld_byte3_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[4] .power_up = "low";

dffeas \W_alu_result[28] (
	.clk(clk_clk),
	.d(\E_alu_result[28]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[28]~q ),
	.prn(vcc));
defparam \W_alu_result[28] .is_wysiwyg = "true";
defparam \W_alu_result[28] .power_up = "low";

dffeas \av_ld_byte3_data[5] (
	.clk(clk_clk),
	.d(src_payload12),
	.asdata(\av_fill_bit~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_aligning_data~q ),
	.ena(!\av_ld_rshift8~0_combout ),
	.q(\av_ld_byte3_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[5] .power_up = "low";

dffeas \W_alu_result[29] (
	.clk(clk_clk),
	.d(\E_alu_result[29]~32_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\W_alu_result[29]~q ),
	.prn(vcc));
defparam \W_alu_result[29] .is_wysiwyg = "true";
defparam \W_alu_result[29] .power_up = "low";

cyclonev_lcell_comb \Add2~85 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[29]~q ),
	.datae(gnd),
	.dataf(!\E_src1[29]~q ),
	.datag(gnd),
	.cin(\Add2~134 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~85_sumout ),
	.cout(\Add2~86 ),
	.shareout());
defparam \Add2~85 .extended_lut = "off";
defparam \Add2~85 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~85 .shared_arith = "off";

cyclonev_lcell_comb \Add2~89 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[25]~q ),
	.datae(gnd),
	.dataf(!\E_src1[25]~q ),
	.datag(gnd),
	.cin(\Add2~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~89_sumout ),
	.cout(\Add2~90 ),
	.shareout());
defparam \Add2~89 .extended_lut = "off";
defparam \Add2~89 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~89 .shared_arith = "off";

cyclonev_lcell_comb \Add2~93 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[27]~q ),
	.datae(gnd),
	.dataf(!\E_src1[27]~q ),
	.datag(gnd),
	.cin(\Add2~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~93_sumout ),
	.cout(\Add2~94 ),
	.shareout());
defparam \Add2~93 .extended_lut = "off";
defparam \Add2~93 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~93 .shared_arith = "off";

cyclonev_lcell_comb \Add2~97 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[19]~q ),
	.datae(gnd),
	.dataf(!\E_src1[19]~q ),
	.datag(gnd),
	.cin(\Add2~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~97_sumout ),
	.cout(\Add2~98 ),
	.shareout());
defparam \Add2~97 .extended_lut = "off";
defparam \Add2~97 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~97 .shared_arith = "off";

cyclonev_lcell_comb \Add2~101 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[20]~q ),
	.datae(gnd),
	.dataf(!\E_src1[20]~q ),
	.datag(gnd),
	.cin(\Add2~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~101_sumout ),
	.cout(\Add2~102 ),
	.shareout());
defparam \Add2~101 .extended_lut = "off";
defparam \Add2~101 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~101 .shared_arith = "off";

cyclonev_lcell_comb \Add2~105 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[21]~q ),
	.datae(gnd),
	.dataf(!\E_src1[21]~q ),
	.datag(gnd),
	.cin(\Add2~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~105_sumout ),
	.cout(\Add2~106 ),
	.shareout());
defparam \Add2~105 .extended_lut = "off";
defparam \Add2~105 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~105 .shared_arith = "off";

cyclonev_lcell_comb \Add2~109 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[22]~q ),
	.datae(gnd),
	.dataf(!\E_src1[22]~q ),
	.datag(gnd),
	.cin(\Add2~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~109_sumout ),
	.cout(\Add2~110 ),
	.shareout());
defparam \Add2~109 .extended_lut = "off";
defparam \Add2~109 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~109 .shared_arith = "off";

cyclonev_lcell_comb \Add2~113 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[23]~q ),
	.datae(gnd),
	.dataf(!\E_src1[23]~q ),
	.datag(gnd),
	.cin(\Add2~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~113_sumout ),
	.cout(\Add2~114 ),
	.shareout());
defparam \Add2~113 .extended_lut = "off";
defparam \Add2~113 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~113 .shared_arith = "off";

cyclonev_lcell_comb \Add2~117 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[24]~q ),
	.datae(gnd),
	.dataf(!\E_src1[24]~q ),
	.datag(gnd),
	.cin(\Add2~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~117_sumout ),
	.cout(\Add2~118 ),
	.shareout());
defparam \Add2~117 .extended_lut = "off";
defparam \Add2~117 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~117 .shared_arith = "off";

cyclonev_lcell_comb \Add2~121 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[18]~q ),
	.datae(gnd),
	.dataf(!\E_src1[18]~q ),
	.datag(gnd),
	.cin(\Add2~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~121_sumout ),
	.cout(\Add2~122 ),
	.shareout());
defparam \Add2~121 .extended_lut = "off";
defparam \Add2~121 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~121 .shared_arith = "off";

cyclonev_lcell_comb \Add2~125 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[17]~q ),
	.datae(gnd),
	.dataf(!\E_src1[17]~q ),
	.datag(gnd),
	.cin(\Add2~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~125_sumout ),
	.cout(\Add2~126 ),
	.shareout());
defparam \Add2~125 .extended_lut = "off";
defparam \Add2~125 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~125 .shared_arith = "off";

cyclonev_lcell_comb \Add2~129 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[26]~q ),
	.datae(gnd),
	.dataf(!\E_src1[26]~q ),
	.datag(gnd),
	.cin(\Add2~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~129_sumout ),
	.cout(\Add2~130 ),
	.shareout());
defparam \Add2~129 .extended_lut = "off";
defparam \Add2~129 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~129 .shared_arith = "off";

cyclonev_lcell_comb \Add2~133 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[28]~q ),
	.datae(gnd),
	.dataf(!\E_src1[28]~q ),
	.datag(gnd),
	.cin(\Add2~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~133_sumout ),
	.cout(\Add2~134 ),
	.shareout());
defparam \Add2~133 .extended_lut = "off";
defparam \Add2~133 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~133 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[6]~9 (
	.dataa(!src0_valid),
	.datab(!\av_ld_byte2_data_nxt[6]~8_combout ),
	.datac(!\av_ld_byte3_data[6]~q ),
	.datad(!q_a_22),
	.datae(!\LessThan0~0_combout ),
	.dataf(!\av_ld_aligning_data~q ),
	.datag(!\av_fill_bit~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[6]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[6]~9 .extended_lut = "on";
defparam \av_ld_byte2_data_nxt[6]~9 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \av_ld_byte2_data_nxt[6]~9 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[5]~13 (
	.dataa(!src0_valid),
	.datab(!\av_ld_byte2_data_nxt[5]~7_combout ),
	.datac(!\av_ld_byte3_data[5]~q ),
	.datad(!q_a_21),
	.datae(!\LessThan0~0_combout ),
	.dataf(!\av_ld_aligning_data~q ),
	.datag(!\av_fill_bit~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[5]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[5]~13 .extended_lut = "on";
defparam \av_ld_byte2_data_nxt[5]~13 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \av_ld_byte2_data_nxt[5]~13 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[4]~17 (
	.dataa(!src0_valid),
	.datab(!\av_ld_byte2_data_nxt[4]~6_combout ),
	.datac(!\av_ld_byte3_data[4]~q ),
	.datad(!q_a_20),
	.datae(!\LessThan0~0_combout ),
	.dataf(!\av_ld_aligning_data~q ),
	.datag(!\av_fill_bit~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[4]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[4]~17 .extended_lut = "on";
defparam \av_ld_byte2_data_nxt[4]~17 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \av_ld_byte2_data_nxt[4]~17 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[1]~21 (
	.dataa(!src0_valid),
	.datab(!\av_ld_byte2_data_nxt[1]~5_combout ),
	.datac(!\av_ld_byte3_data[1]~q ),
	.datad(!q_a_17),
	.datae(!\LessThan0~0_combout ),
	.dataf(!\av_ld_aligning_data~q ),
	.datag(!\av_fill_bit~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[1]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[1]~21 .extended_lut = "on";
defparam \av_ld_byte2_data_nxt[1]~21 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \av_ld_byte2_data_nxt[1]~21 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[2]~25 (
	.dataa(!src0_valid),
	.datab(!\av_ld_byte2_data_nxt[2]~4_combout ),
	.datac(!\av_ld_byte3_data[2]~q ),
	.datad(!q_a_18),
	.datae(!\LessThan0~0_combout ),
	.dataf(!\av_ld_aligning_data~q ),
	.datag(!\av_fill_bit~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[2]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[2]~25 .extended_lut = "on";
defparam \av_ld_byte2_data_nxt[2]~25 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \av_ld_byte2_data_nxt[2]~25 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[3]~29 (
	.dataa(!src0_valid),
	.datab(!\av_ld_byte2_data_nxt[3]~3_combout ),
	.datac(!\av_ld_byte3_data[3]~q ),
	.datad(!q_a_19),
	.datae(!\LessThan0~0_combout ),
	.dataf(!\av_ld_aligning_data~q ),
	.datag(!\av_fill_bit~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[3]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[3]~29 .extended_lut = "on";
defparam \av_ld_byte2_data_nxt[3]~29 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \av_ld_byte2_data_nxt[3]~29 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[0]~33 (
	.dataa(!src0_valid),
	.datab(!\av_ld_byte2_data_nxt[0]~2_combout ),
	.datac(!\av_ld_byte3_data[0]~q ),
	.datad(!q_a_16),
	.datae(!\LessThan0~0_combout ),
	.dataf(!\av_ld_aligning_data~q ),
	.datag(!\av_fill_bit~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[0]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[0]~33 .extended_lut = "on";
defparam \av_ld_byte2_data_nxt[0]~33 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \av_ld_byte2_data_nxt[0]~33 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[7]~9 (
	.dataa(!src0_valid),
	.datab(!\av_ld_byte1_data_nxt[7]~8_combout ),
	.datac(!\av_ld_byte2_data[7]~q ),
	.datad(!q_a_15),
	.datae(!\LessThan0~0_combout ),
	.dataf(!\av_ld_aligning_data~q ),
	.datag(!\av_fill_bit~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[7]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[7]~9 .extended_lut = "on";
defparam \av_ld_byte1_data_nxt[7]~9 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \av_ld_byte1_data_nxt[7]~9 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[6]~13 (
	.dataa(!src0_valid),
	.datab(!\av_ld_byte1_data_nxt[6]~7_combout ),
	.datac(!\av_ld_byte2_data[6]~q ),
	.datad(!q_a_14),
	.datae(!\LessThan0~0_combout ),
	.dataf(!\av_ld_aligning_data~q ),
	.datag(!\av_fill_bit~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[6]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[6]~13 .extended_lut = "on";
defparam \av_ld_byte1_data_nxt[6]~13 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \av_ld_byte1_data_nxt[6]~13 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[5]~17 (
	.dataa(!src0_valid),
	.datab(!\av_ld_byte1_data_nxt[5]~6_combout ),
	.datac(!\av_ld_byte2_data[5]~q ),
	.datad(!q_a_13),
	.datae(!\LessThan0~0_combout ),
	.dataf(!\av_ld_aligning_data~q ),
	.datag(!\av_fill_bit~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[5]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[5]~17 .extended_lut = "on";
defparam \av_ld_byte1_data_nxt[5]~17 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \av_ld_byte1_data_nxt[5]~17 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[4]~21 (
	.dataa(!src0_valid),
	.datab(!\av_ld_byte1_data_nxt[4]~5_combout ),
	.datac(!\av_ld_byte2_data[4]~q ),
	.datad(!q_a_12),
	.datae(!\LessThan0~0_combout ),
	.dataf(!\av_ld_aligning_data~q ),
	.datag(!\av_fill_bit~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[4]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[4]~21 .extended_lut = "on";
defparam \av_ld_byte1_data_nxt[4]~21 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \av_ld_byte1_data_nxt[4]~21 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[1]~25 (
	.dataa(!src0_valid),
	.datab(!\av_ld_byte1_data_nxt[1]~4_combout ),
	.datac(!\av_ld_byte2_data[1]~q ),
	.datad(!q_a_9),
	.datae(!\LessThan0~0_combout ),
	.dataf(!\av_ld_aligning_data~q ),
	.datag(!\av_fill_bit~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[1]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[1]~25 .extended_lut = "on";
defparam \av_ld_byte1_data_nxt[1]~25 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \av_ld_byte1_data_nxt[1]~25 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[2]~29 (
	.dataa(!src0_valid),
	.datab(!\av_ld_byte1_data_nxt[2]~3_combout ),
	.datac(!\av_ld_byte2_data[2]~q ),
	.datad(!q_a_10),
	.datae(!\LessThan0~0_combout ),
	.dataf(!\av_ld_aligning_data~q ),
	.datag(!\av_fill_bit~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[2]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[2]~29 .extended_lut = "on";
defparam \av_ld_byte1_data_nxt[2]~29 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \av_ld_byte1_data_nxt[2]~29 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[0]~33 (
	.dataa(!src0_valid),
	.datab(!\av_ld_byte1_data_nxt[0]~2_combout ),
	.datac(!\av_ld_byte2_data[0]~q ),
	.datad(!q_a_8),
	.datae(!\LessThan0~0_combout ),
	.dataf(!\av_ld_aligning_data~q ),
	.datag(!\av_fill_bit~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[0]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[0]~33 .extended_lut = "on";
defparam \av_ld_byte1_data_nxt[0]~33 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \av_ld_byte1_data_nxt[0]~33 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[0]~31 (
	.dataa(!\W_cmp_result~q ),
	.datab(!\av_ld_byte0_data[0]~q ),
	.datac(!\W_control_rd_data[0]~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\R_ctrl_rd_ctl_reg~q ),
	.dataf(!\R_ctrl_br_cmp~q ),
	.datag(!\W_alu_result[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[0]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[0]~31 .extended_lut = "on";
defparam \W_rf_wr_data[0]~31 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \W_rf_wr_data[0]~31 .shared_arith = "off";

dffeas R_wr_dst_reg(
	.clk(clk_clk),
	.d(\D_wr_dst_reg~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_wr_dst_reg~q ),
	.prn(vcc));
defparam R_wr_dst_reg.is_wysiwyg = "true";
defparam R_wr_dst_reg.power_up = "low";

cyclonev_lcell_comb W_rf_wren(
	.dataa(!r_sync_rst),
	.datab(!\R_wr_dst_reg~q ),
	.datac(!\W_valid~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wren~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam W_rf_wren.extended_lut = "off";
defparam W_rf_wren.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam W_rf_wren.shared_arith = "off";

dffeas \W_control_rd_data[0] (
	.clk(clk_clk),
	.d(\E_control_rd_data[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_control_rd_data[0]~q ),
	.prn(vcc));
defparam \W_control_rd_data[0] .is_wysiwyg = "true";
defparam \W_control_rd_data[0] .power_up = "low";

dffeas \R_dst_regnum[0] (
	.clk(clk_clk),
	.d(\D_dst_regnum[0]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[0]~q ),
	.prn(vcc));
defparam \R_dst_regnum[0] .is_wysiwyg = "true";
defparam \R_dst_regnum[0] .power_up = "low";

dffeas \R_dst_regnum[1] (
	.clk(clk_clk),
	.d(\D_dst_regnum[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[1]~q ),
	.prn(vcc));
defparam \R_dst_regnum[1] .is_wysiwyg = "true";
defparam \R_dst_regnum[1] .power_up = "low";

dffeas \R_dst_regnum[2] (
	.clk(clk_clk),
	.d(\D_dst_regnum[2]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[2]~q ),
	.prn(vcc));
defparam \R_dst_regnum[2] .is_wysiwyg = "true";
defparam \R_dst_regnum[2] .power_up = "low";

dffeas \R_dst_regnum[3] (
	.clk(clk_clk),
	.d(\D_dst_regnum[3]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[3]~q ),
	.prn(vcc));
defparam \R_dst_regnum[3] .is_wysiwyg = "true";
defparam \R_dst_regnum[3] .power_up = "low";

dffeas \R_dst_regnum[4] (
	.clk(clk_clk),
	.d(\D_dst_regnum[4]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[4]~q ),
	.prn(vcc));
defparam \R_dst_regnum[4] .is_wysiwyg = "true";
defparam \R_dst_regnum[4] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[1]~0 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte0_data[1]~q ),
	.datae(!\W_alu_result[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[1]~0 .extended_lut = "off";
defparam \W_rf_wr_data[1]~0 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[2]~1 (
	.dataa(!W_alu_result_2),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte0_data[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[2]~1 .extended_lut = "off";
defparam \W_rf_wr_data[2]~1 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[3]~2 (
	.dataa(!W_alu_result_3),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte0_data[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[3]~2 .extended_lut = "off";
defparam \W_rf_wr_data[3]~2 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[4]~3 (
	.dataa(!W_alu_result_4),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte0_data[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[4]~3 .extended_lut = "off";
defparam \W_rf_wr_data[4]~3 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[4]~3 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[5]~4 (
	.dataa(!W_alu_result_5),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte0_data[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[5]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[5]~4 .extended_lut = "off";
defparam \W_rf_wr_data[5]~4 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[5]~4 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[1]~0 (
	.dataa(!\D_iw[23]~q ),
	.datab(!\D_iw[18]~q ),
	.datac(!\D_ctrl_b_is_dst~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[1]~0 .extended_lut = "off";
defparam \D_dst_regnum[1]~0 .lut_mask = 64'h5353535353535353;
defparam \D_dst_regnum[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[1]~1 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal0~7_combout ),
	.datac(!\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.datad(!\D_ctrl_implicit_dst_eretaddr~1_combout ),
	.datae(!\D_ctrl_exception~0_combout ),
	.dataf(!\D_dst_regnum[1]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[1]~1 .extended_lut = "off";
defparam \D_dst_regnum[1]~1 .lut_mask = 64'hFFFBFFFFFFFFFFFF;
defparam \D_dst_regnum[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[2]~2 (
	.dataa(!\D_iw[24]~q ),
	.datab(!\D_iw[19]~q ),
	.datac(!\D_ctrl_b_is_dst~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[2]~2 .extended_lut = "off";
defparam \D_dst_regnum[2]~2 .lut_mask = 64'h5353535353535353;
defparam \D_dst_regnum[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[2]~3 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal0~7_combout ),
	.datac(!\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.datad(!\D_ctrl_implicit_dst_eretaddr~1_combout ),
	.datae(!\D_ctrl_exception~0_combout ),
	.dataf(!\D_dst_regnum[2]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[2]~3 .extended_lut = "off";
defparam \D_dst_regnum[2]~3 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \D_dst_regnum[2]~3 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[0]~4 (
	.dataa(!\D_iw[22]~q ),
	.datab(!\D_iw[17]~q ),
	.datac(!\D_ctrl_b_is_dst~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[0]~4 .extended_lut = "off";
defparam \D_dst_regnum[0]~4 .lut_mask = 64'h5353535353535353;
defparam \D_dst_regnum[0]~4 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[0]~5 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal0~7_combout ),
	.datac(!\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.datad(!\D_ctrl_implicit_dst_eretaddr~1_combout ),
	.datae(!\D_ctrl_exception~0_combout ),
	.dataf(!\D_dst_regnum[0]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[0]~5 .extended_lut = "off";
defparam \D_dst_regnum[0]~5 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \D_dst_regnum[0]~5 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[3]~6 (
	.dataa(!\D_iw[25]~q ),
	.datab(!\D_iw[20]~q ),
	.datac(!\D_ctrl_b_is_dst~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[3]~6 .extended_lut = "off";
defparam \D_dst_regnum[3]~6 .lut_mask = 64'h5353535353535353;
defparam \D_dst_regnum[3]~6 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[3]~7 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal0~7_combout ),
	.datac(!\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.datad(!\D_ctrl_implicit_dst_eretaddr~1_combout ),
	.datae(!\D_ctrl_exception~0_combout ),
	.dataf(!\D_dst_regnum[3]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[3]~7 .extended_lut = "off";
defparam \D_dst_regnum[3]~7 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \D_dst_regnum[3]~7 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[4]~8 (
	.dataa(!\D_iw[26]~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\D_ctrl_b_is_dst~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[4]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[4]~8 .extended_lut = "off";
defparam \D_dst_regnum[4]~8 .lut_mask = 64'h5353535353535353;
defparam \D_dst_regnum[4]~8 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[4]~9 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal0~7_combout ),
	.datac(!\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.datad(!\D_ctrl_implicit_dst_eretaddr~1_combout ),
	.datae(!\D_ctrl_exception~0_combout ),
	.dataf(!\D_dst_regnum[4]~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[4]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[4]~9 .extended_lut = "off";
defparam \D_dst_regnum[4]~9 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \D_dst_regnum[4]~9 .shared_arith = "off";

cyclonev_lcell_comb \D_wr_dst_reg~0 (
	.dataa(!\Equal0~11_combout ),
	.datab(!\R_ctrl_br_nxt~2_combout ),
	.datac(!\R_src2_use_imm~5_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_wr_dst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_wr_dst_reg~0 .extended_lut = "off";
defparam \D_wr_dst_reg~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \D_wr_dst_reg~0 .shared_arith = "off";

cyclonev_lcell_comb D_wr_dst_reg(
	.dataa(!\D_dst_regnum[1]~1_combout ),
	.datab(!\D_dst_regnum[2]~3_combout ),
	.datac(!\D_dst_regnum[0]~5_combout ),
	.datad(!\D_dst_regnum[3]~7_combout ),
	.datae(!\D_dst_regnum[4]~9_combout ),
	.dataf(!\D_wr_dst_reg~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_wr_dst_reg~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_wr_dst_reg.extended_lut = "off";
defparam D_wr_dst_reg.lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam D_wr_dst_reg.shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_ld_signed~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[4]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_ld_signed~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_ld_signed~0 .extended_lut = "off";
defparam \D_ctrl_ld_signed~0 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \D_ctrl_ld_signed~0 .shared_arith = "off";

dffeas \av_ld_byte1_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data_nxt[0]~33_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[0] .power_up = "low";

cyclonev_lcell_comb \av_ld_rshift8~0 (
	.dataa(!\W_alu_result[0]~q ),
	.datab(!\W_alu_result[1]~q ),
	.datac(!\av_ld_aligning_data~q ),
	.datad(!\av_ld_align_cycle[1]~q ),
	.datae(!\av_ld_align_cycle[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_rshift8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_rshift8~0 .extended_lut = "off";
defparam \av_ld_rshift8~0 .lut_mask = 64'hFFFFFF7FFFFFFF7F;
defparam \av_ld_rshift8~0 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte0_data[2]~0 (
	.dataa(!\W_alu_result[0]~q ),
	.datab(!\W_alu_result[1]~q ),
	.datac(!\av_ld_aligning_data~q ),
	.datad(!\av_ld_align_cycle[1]~q ),
	.datae(!\av_ld_align_cycle[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte0_data[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte0_data[2]~0 .extended_lut = "off";
defparam \av_ld_byte0_data[2]~0 .lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam \av_ld_byte0_data[2]~0 .shared_arith = "off";

dffeas W_status_reg_pie(
	.clk(clk_clk),
	.d(\W_status_reg_pie_inst_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_status_reg_pie~q ),
	.prn(vcc));
defparam W_status_reg_pie.is_wysiwyg = "true";
defparam W_status_reg_pie.power_up = "low";

cyclonev_lcell_comb \Equal133~0 (
	.dataa(!\D_iw[8]~q ),
	.datab(!\D_iw[10]~q ),
	.datac(!\D_iw[9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal133~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal133~0 .extended_lut = "off";
defparam \Equal133~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \Equal133~0 .shared_arith = "off";

dffeas W_bstatus_reg(
	.clk(clk_clk),
	.d(\W_bstatus_reg_inst_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_bstatus_reg~q ),
	.prn(vcc));
defparam W_bstatus_reg.is_wysiwyg = "true";
defparam W_bstatus_reg.power_up = "low";

cyclonev_lcell_comb \E_control_rd_data[0]~0 (
	.dataa(!\D_iw[6]~q ),
	.datab(!\D_iw[7]~q ),
	.datac(!\W_status_reg_pie~q ),
	.datad(!\Equal133~0_combout ),
	.datae(!\W_estatus_reg~q ),
	.dataf(!\W_bstatus_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_control_rd_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_control_rd_data[0]~0 .extended_lut = "off";
defparam \E_control_rd_data[0]~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \E_control_rd_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[0]~16 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_logic_result[0]~23_combout ),
	.datad(!\E_shift_rot_result[0]~q ),
	.datae(!\Add2~69_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[0]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[0]~16 .extended_lut = "off";
defparam \E_alu_result[0]~16 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[0]~16 .shared_arith = "off";

dffeas \av_ld_byte1_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data_nxt[3]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[3] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[11]~5 (
	.dataa(!W_alu_result_11),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte1_data[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[11]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[11]~5 .extended_lut = "off";
defparam \W_rf_wr_data[11]~5 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[11]~5 .shared_arith = "off";

dffeas \av_ld_byte1_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data_nxt[2]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[2] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[10]~6 (
	.dataa(!W_alu_result_10),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte1_data[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[10]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[10]~6 .extended_lut = "off";
defparam \W_rf_wr_data[10]~6 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[10]~6 .shared_arith = "off";

dffeas \av_ld_byte1_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data_nxt[1]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[1] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[9]~7 (
	.dataa(!W_alu_result_9),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte1_data[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[9]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[9]~7 .extended_lut = "off";
defparam \W_rf_wr_data[9]~7 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[9]~7 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[8]~8 (
	.dataa(!W_alu_result_8),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte1_data[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[8]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[8]~8 .extended_lut = "off";
defparam \W_rf_wr_data[8]~8 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[8]~8 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[7]~9 (
	.dataa(!W_alu_result_7),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte0_data[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[7]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[7]~9 .extended_lut = "off";
defparam \W_rf_wr_data[7]~9 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[7]~9 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[6]~10 (
	.dataa(!W_alu_result_6),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte0_data[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[6]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[6]~10 .extended_lut = "off";
defparam \W_rf_wr_data[6]~10 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[6]~10 .shared_arith = "off";

dffeas \av_ld_byte1_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data_nxt[4]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[4] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[12]~11 (
	.dataa(!W_alu_result_12),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte1_data[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[12]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[12]~11 .extended_lut = "off";
defparam \W_rf_wr_data[12]~11 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[12]~11 .shared_arith = "off";

dffeas \av_ld_byte1_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data_nxt[5]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[5] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[13]~12 (
	.dataa(!W_alu_result_13),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte1_data[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[13]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[13]~12 .extended_lut = "off";
defparam \W_rf_wr_data[13]~12 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[13]~12 .shared_arith = "off";

dffeas \av_ld_byte1_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data_nxt[6]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[6] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[14]~13 (
	.dataa(!W_alu_result_14),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte1_data[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[14]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[14]~13 .extended_lut = "off";
defparam \W_rf_wr_data[14]~13 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[14]~13 .shared_arith = "off";

dffeas \av_ld_byte1_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data_nxt[7]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[7] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[15]~14 (
	.dataa(!W_alu_result_15),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte1_data[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[15]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[15]~14 .extended_lut = "off";
defparam \W_rf_wr_data[15]~14 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[15]~14 .shared_arith = "off";

dffeas \av_ld_byte2_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data_nxt[0]~33_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_byte2_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[0] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[16]~15 (
	.dataa(!W_alu_result_16),
	.datab(!\R_ctrl_rd_ctl_reg~q ),
	.datac(!\R_ctrl_br_cmp~q ),
	.datad(!\R_ctrl_ld~q ),
	.datae(!\av_ld_byte2_data[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[16]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[16]~15 .extended_lut = "off";
defparam \W_rf_wr_data[16]~15 .lut_mask = 64'hDDF5FFFFDDF5FFFF;
defparam \W_rf_wr_data[16]~15 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[1]~26 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[1]~q ),
	.datad(!\E_src1[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[1]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[1]~26 .extended_lut = "off";
defparam \E_logic_result[1]~26 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[1]~26 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[1]~17 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[1]~q ),
	.datad(!\Add2~61_sumout ),
	.datae(!\E_logic_result[1]~26_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[1]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[1]~17 .extended_lut = "off";
defparam \E_alu_result[1]~17 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[1]~17 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\W_alu_result[0]~q ),
	.datab(!\W_alu_result[1]~q ),
	.datac(!\av_ld_align_cycle[1]~q ),
	.datad(!\av_ld_align_cycle[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \LessThan0~0 .shared_arith = "off";

dffeas R_ctrl_ld_signed(
	.clk(clk_clk),
	.d(\D_ctrl_ld_signed~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_ld_signed~q ),
	.prn(vcc));
defparam R_ctrl_ld_signed.is_wysiwyg = "true";
defparam R_ctrl_ld_signed.power_up = "low";

cyclonev_lcell_comb \av_fill_bit~0 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_ctrl_mem16~0_combout ),
	.datac(!\av_ld_byte0_data[7]~q ),
	.datad(!\av_ld_byte1_data[7]~q ),
	.datae(!\R_ctrl_ld_signed~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_fill_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_fill_bit~0 .extended_lut = "off";
defparam \av_fill_bit~0 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \av_fill_bit~0 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_en~0 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_ctrl_mem16~0_combout ),
	.datac(!\av_ld_byte0_data[2]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_en~0 .extended_lut = "off";
defparam \av_ld_byte1_data_en~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \av_ld_byte1_data_en~0 .shared_arith = "off";

dffeas R_ctrl_wrctl_inst(
	.clk(clk_clk),
	.d(\D_op_wrctl~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_wrctl_inst~q ),
	.prn(vcc));
defparam R_ctrl_wrctl_inst.is_wysiwyg = "true";
defparam R_ctrl_wrctl_inst.power_up = "low";

cyclonev_lcell_comb \W_status_reg_pie_inst_nxt~0 (
	.dataa(!\D_iw[8]~q ),
	.datab(!\D_iw[10]~q ),
	.datac(!\D_iw[9]~q ),
	.datad(!\D_iw[6]~q ),
	.datae(!\D_iw[7]~q ),
	.dataf(!\R_ctrl_wrctl_inst~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_status_reg_pie_inst_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_status_reg_pie_inst_nxt~0 .extended_lut = "off";
defparam \W_status_reg_pie_inst_nxt~0 .lut_mask = 64'hFFFFFFFEFFFFFFFF;
defparam \W_status_reg_pie_inst_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \W_status_reg_pie_inst_nxt~1 (
	.dataa(!\E_src1[0]~q ),
	.datab(!\Equal0~0_combout ),
	.datac(!\W_status_reg_pie~q ),
	.datad(!\W_bstatus_reg~q ),
	.datae(!\Equal62~16_combout ),
	.dataf(!\W_status_reg_pie_inst_nxt~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_status_reg_pie_inst_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_status_reg_pie_inst_nxt~1 .extended_lut = "off";
defparam \W_status_reg_pie_inst_nxt~1 .lut_mask = 64'hDFFF7FFF7FFFDFFF;
defparam \W_status_reg_pie_inst_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \W_status_reg_pie_inst_nxt~2 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\W_estatus_reg~q ),
	.datac(!\Equal62~15_combout ),
	.datad(!\R_ctrl_exception~q ),
	.datae(!\R_ctrl_break~q ),
	.dataf(!\W_status_reg_pie_inst_nxt~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_status_reg_pie_inst_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_status_reg_pie_inst_nxt~2 .extended_lut = "off";
defparam \W_status_reg_pie_inst_nxt~2 .lut_mask = 64'hFFFFFF7BFFFFFFFF;
defparam \W_status_reg_pie_inst_nxt~2 .shared_arith = "off";

cyclonev_lcell_comb \W_estatus_reg_inst_nxt~0 (
	.dataa(!\E_src1[0]~q ),
	.datab(!\D_iw[6]~q ),
	.datac(!\D_iw[7]~q ),
	.datad(!\Equal133~0_combout ),
	.datae(!\W_estatus_reg~q ),
	.dataf(!\R_ctrl_wrctl_inst~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_estatus_reg_inst_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_estatus_reg_inst_nxt~0 .extended_lut = "off";
defparam \W_estatus_reg_inst_nxt~0 .lut_mask = 64'h7DD7FFFFD77DFFFF;
defparam \W_estatus_reg_inst_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \E_wrctl_bstatus~0 (
	.dataa(!\D_iw[6]~q ),
	.datab(!\D_iw[7]~q ),
	.datac(!\Equal133~0_combout ),
	.datad(!\R_ctrl_wrctl_inst~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_wrctl_bstatus~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_wrctl_bstatus~0 .extended_lut = "off";
defparam \E_wrctl_bstatus~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \E_wrctl_bstatus~0 .shared_arith = "off";

cyclonev_lcell_comb \W_bstatus_reg_inst_nxt~0 (
	.dataa(!\E_src1[0]~q ),
	.datab(!\W_status_reg_pie~q ),
	.datac(!\W_bstatus_reg~q ),
	.datad(!\R_ctrl_break~q ),
	.datae(!\E_wrctl_bstatus~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_bstatus_reg_inst_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_bstatus_reg_inst_nxt~0 .extended_lut = "off";
defparam \W_bstatus_reg_inst_nxt~0 .lut_mask = 64'h7FFFFF7F7FFFFF7F;
defparam \W_bstatus_reg_inst_nxt~0 .shared_arith = "off";

dffeas \av_ld_byte2_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data_nxt[3]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_byte2_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[3] .power_up = "low";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[3]~0 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\LessThan0~0_combout ),
	.datac(!\av_fill_bit~0_combout ),
	.datad(!src0_valid),
	.datae(!q_a_11),
	.dataf(!\av_ld_byte1_data_nxt[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[3]~0 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[3]~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \av_ld_byte1_data_nxt[3]~0 .shared_arith = "off";

dffeas \av_ld_byte2_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data_nxt[2]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_byte2_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[2] .power_up = "low";

dffeas \av_ld_byte2_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data_nxt[1]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_byte2_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[1] .power_up = "low";

dffeas \av_ld_byte2_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data_nxt[4]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_byte2_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[4] .power_up = "low";

dffeas \av_ld_byte2_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data_nxt[5]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_byte2_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[5] .power_up = "low";

dffeas \av_ld_byte2_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data_nxt[6]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_byte2_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[6] .power_up = "low";

dffeas \av_ld_byte2_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data_nxt[7]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_byte2_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[7] .power_up = "low";

cyclonev_lcell_comb \W_rf_wr_data[25]~16 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte3_data[1]~q ),
	.datae(!\W_alu_result[25]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[25]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[25]~16 .extended_lut = "off";
defparam \W_rf_wr_data[25]~16 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[25]~16 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[27]~17 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte3_data[3]~q ),
	.datae(!\W_alu_result[27]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[27]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[27]~17 .extended_lut = "off";
defparam \W_rf_wr_data[27]~17 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[27]~17 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[19]~18 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte2_data[3]~q ),
	.datae(!\W_alu_result[19]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[19]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[19]~18 .extended_lut = "off";
defparam \W_rf_wr_data[19]~18 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[19]~18 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[20]~19 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte2_data[4]~q ),
	.datae(!\W_alu_result[20]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[20]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[20]~19 .extended_lut = "off";
defparam \W_rf_wr_data[20]~19 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[20]~19 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[21]~20 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte2_data[5]~q ),
	.datae(!\W_alu_result[21]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[21]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[21]~20 .extended_lut = "off";
defparam \W_rf_wr_data[21]~20 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[21]~20 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[22]~21 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte2_data[6]~q ),
	.datae(!\W_alu_result[22]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[22]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[22]~21 .extended_lut = "off";
defparam \W_rf_wr_data[22]~21 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[22]~21 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[23]~22 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte2_data[7]~q ),
	.datae(!\W_alu_result[23]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[23]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[23]~22 .extended_lut = "off";
defparam \W_rf_wr_data[23]~22 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[23]~22 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[24]~23 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte3_data[0]~q ),
	.datae(!\W_alu_result[24]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[24]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[24]~23 .extended_lut = "off";
defparam \W_rf_wr_data[24]~23 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[24]~23 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[18]~24 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte2_data[2]~q ),
	.datae(!\W_alu_result[18]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[18]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[18]~24 .extended_lut = "off";
defparam \W_rf_wr_data[18]~24 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[18]~24 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[17]~25 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte2_data[1]~q ),
	.datae(!\W_alu_result[17]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[17]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[17]~25 .extended_lut = "off";
defparam \W_rf_wr_data[17]~25 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[17]~25 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[26]~26 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte3_data[2]~q ),
	.datae(!\W_alu_result[26]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[26]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[26]~26 .extended_lut = "off";
defparam \W_rf_wr_data[26]~26 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[26]~26 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[31]~27 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte3_data[7]~q ),
	.datae(!\W_alu_result[31]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[31]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[31]~27 .extended_lut = "off";
defparam \W_rf_wr_data[31]~27 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[31]~27 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[30]~28 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte3_data[6]~q ),
	.datae(!\W_alu_result[30]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[30]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[30]~28 .extended_lut = "off";
defparam \W_rf_wr_data[30]~28 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[30]~28 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[28]~29 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte3_data[4]~q ),
	.datae(!\W_alu_result[28]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[28]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[28]~29 .extended_lut = "off";
defparam \W_rf_wr_data[28]~29 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[28]~29 .shared_arith = "off";

cyclonev_lcell_comb \W_rf_wr_data[29]~30 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\av_ld_byte3_data[5]~q ),
	.datae(!\W_alu_result[29]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_rf_wr_data[29]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_rf_wr_data[29]~30 .extended_lut = "off";
defparam \W_rf_wr_data[29]~30 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \W_rf_wr_data[29]~30 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~17 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~17 .extended_lut = "off";
defparam \Equal62~17 .lut_mask = 64'hFFFFBFFFFFFFFFFF;
defparam \Equal62~17 .shared_arith = "off";

cyclonev_lcell_comb D_op_wrctl(
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal62~17_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_op_wrctl~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_op_wrctl.extended_lut = "off";
defparam D_op_wrctl.lut_mask = 64'h7777777777777777;
defparam D_op_wrctl.shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[7]~0 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\LessThan0~0_combout ),
	.datac(!\av_fill_bit~0_combout ),
	.datad(!src0_valid),
	.datae(!q_a_23),
	.dataf(!\av_ld_byte2_data_nxt[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[7]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[7]~0 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[7]~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \av_ld_byte2_data_nxt[7]~0 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[25]~18 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_logic_result[25]~15_combout ),
	.datad(!\E_shift_rot_result[25]~q ),
	.datae(!\Add2~89_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[25]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[25]~18 .extended_lut = "off";
defparam \E_alu_result[25]~18 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[25]~18 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[27]~19 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_logic_result[27]~16_combout ),
	.datad(!\E_shift_rot_result[27]~q ),
	.datae(!\Add2~93_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[27]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[27]~19 .extended_lut = "off";
defparam \E_alu_result[27]~19 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[27]~19 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[19]~20 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_logic_result[19]~17_combout ),
	.datad(!\E_shift_rot_result[19]~q ),
	.datae(!\Add2~97_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[19]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[19]~20 .extended_lut = "off";
defparam \E_alu_result[19]~20 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[19]~20 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[20]~21 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_logic_result[20]~18_combout ),
	.datad(!\E_shift_rot_result[20]~q ),
	.datae(!\Add2~101_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[20]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[20]~21 .extended_lut = "off";
defparam \E_alu_result[20]~21 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[20]~21 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[21]~22 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_logic_result[21]~19_combout ),
	.datad(!\E_shift_rot_result[21]~q ),
	.datae(!\Add2~105_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[21]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[21]~22 .extended_lut = "off";
defparam \E_alu_result[21]~22 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[21]~22 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[22]~23 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_logic_result[22]~20_combout ),
	.datad(!\E_shift_rot_result[22]~q ),
	.datae(!\Add2~109_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[22]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[22]~23 .extended_lut = "off";
defparam \E_alu_result[22]~23 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[22]~23 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[23]~24 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_logic_result[23]~21_combout ),
	.datad(!\E_shift_rot_result[23]~q ),
	.datae(!\Add2~113_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[23]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[23]~24 .extended_lut = "off";
defparam \E_alu_result[23]~24 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[23]~24 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[24]~25 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_logic_result[24]~22_combout ),
	.datad(!\E_shift_rot_result[24]~q ),
	.datae(!\Add2~117_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[24]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[24]~25 .extended_lut = "off";
defparam \E_alu_result[24]~25 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[24]~25 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[18]~27 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[18]~q ),
	.datad(!\E_src1[18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[18]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[18]~27 .extended_lut = "off";
defparam \E_logic_result[18]~27 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[18]~27 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[18]~26 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_logic_result[18]~27_combout ),
	.datad(!\E_shift_rot_result[18]~q ),
	.datae(!\Add2~121_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[18]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[18]~26 .extended_lut = "off";
defparam \E_alu_result[18]~26 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[18]~26 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[17]~28 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[17]~q ),
	.datad(!\E_src1[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[17]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[17]~28 .extended_lut = "off";
defparam \E_logic_result[17]~28 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[17]~28 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[17]~27 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[17]~q ),
	.datad(!\E_logic_result[17]~28_combout ),
	.datae(!\Add2~125_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[17]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[17]~27 .extended_lut = "off";
defparam \E_alu_result[17]~27 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[17]~27 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[26]~29 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[26]~q ),
	.datad(!\E_src1[26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[26]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[26]~29 .extended_lut = "off";
defparam \E_logic_result[26]~29 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[26]~29 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[26]~28 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_logic_result[26]~29_combout ),
	.datad(!\E_shift_rot_result[26]~q ),
	.datae(!\Add2~129_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[26]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[26]~28 .extended_lut = "off";
defparam \E_alu_result[26]~28 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[26]~28 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[31]~30 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[31]~q ),
	.datad(!\E_src1[31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[31]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[31]~30 .extended_lut = "off";
defparam \E_logic_result[31]~30 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[31]~30 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[31]~29 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_logic_result[31]~30_combout ),
	.datad(!\Add2~73_sumout ),
	.datae(!\E_shift_rot_result[31]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[31]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[31]~29 .extended_lut = "off";
defparam \E_alu_result[31]~29 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[31]~29 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[30]~31 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[30]~q ),
	.datad(!\E_src1[30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[30]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[30]~31 .extended_lut = "off";
defparam \E_logic_result[30]~31 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[30]~31 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[30]~30 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_logic_result[30]~31_combout ),
	.datad(!\Add2~81_sumout ),
	.datae(!\E_shift_rot_result[30]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[30]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[30]~30 .extended_lut = "off";
defparam \E_alu_result[30]~30 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[30]~30 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[28]~31 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_logic_result[28]~24_combout ),
	.datad(!\E_shift_rot_result[28]~q ),
	.datae(!\Add2~133_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[28]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[28]~31 .extended_lut = "off";
defparam \E_alu_result[28]~31 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[28]~31 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[29]~32 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_logic_result[29]~25_combout ),
	.datad(!\Add2~85_sumout ),
	.datae(!\E_shift_rot_result[29]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[29]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[29]~32 .extended_lut = "off";
defparam \E_alu_result[29]~32 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[29]~32 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[3]~1 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\av_ld_byte2_data[3]~q ),
	.datac(!src0_valid1),
	.datad(!av_readdata_pre_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[3]~1 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[3]~1 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \av_ld_byte1_data_nxt[3]~1 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[7]~1 (
	.dataa(!\av_ld_aligning_data~q ),
	.datab(!\av_ld_byte3_data[7]~q ),
	.datac(!src0_valid1),
	.datad(!av_readdata_pre_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[7]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[7]~1 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[7]~1 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \av_ld_byte2_data_nxt[7]~1 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[0]~2 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_8),
	.datad(!av_readdata_pre_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[0]~2 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[0]~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \av_ld_byte1_data_nxt[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[2]~3 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_10),
	.datad(!av_readdata_pre_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[2]~3 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[2]~3 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \av_ld_byte1_data_nxt[2]~3 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[1]~4 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_9),
	.datad(!av_readdata_pre_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[1]~4 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[1]~4 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \av_ld_byte1_data_nxt[1]~4 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[4]~5 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_12),
	.datad(!av_readdata_pre_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[4]~5 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[4]~5 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \av_ld_byte1_data_nxt[4]~5 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[5]~6 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_13),
	.datad(!av_readdata_pre_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[5]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[5]~6 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[5]~6 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \av_ld_byte1_data_nxt[5]~6 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[6]~7 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_14),
	.datad(!av_readdata_pre_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[6]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[6]~7 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[6]~7 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \av_ld_byte1_data_nxt[6]~7 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data_nxt[7]~8 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_15),
	.datad(!av_readdata_pre_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data_nxt[7]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data_nxt[7]~8 .extended_lut = "off";
defparam \av_ld_byte1_data_nxt[7]~8 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \av_ld_byte1_data_nxt[7]~8 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[0]~2 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_161),
	.datad(!av_readdata_pre_16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[0]~2 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[0]~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \av_ld_byte2_data_nxt[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[3]~3 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_191),
	.datad(!av_readdata_pre_19),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[3]~3 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[3]~3 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \av_ld_byte2_data_nxt[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[2]~4 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_181),
	.datad(!av_readdata_pre_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[2]~4 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[2]~4 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \av_ld_byte2_data_nxt[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[1]~5 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_171),
	.datad(!av_readdata_pre_17),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[1]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[1]~5 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[1]~5 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \av_ld_byte2_data_nxt[1]~5 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[4]~6 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_201),
	.datad(!av_readdata_pre_20),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[4]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[4]~6 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[4]~6 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \av_ld_byte2_data_nxt[4]~6 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[5]~7 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_211),
	.datad(!av_readdata_pre_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[5]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[5]~7 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[5]~7 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \av_ld_byte2_data_nxt[5]~7 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte2_data_nxt[6]~8 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_221),
	.datad(!av_readdata_pre_22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte2_data_nxt[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte2_data_nxt[6]~8 .extended_lut = "off";
defparam \av_ld_byte2_data_nxt[6]~8 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \av_ld_byte2_data_nxt[6]~8 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_implicit_dst_eretaddr~1 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\D_iw[12]~q ),
	.datad(!\D_iw[11]~q ),
	.datae(!\D_iw[16]~q ),
	.dataf(!\D_iw[15]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_implicit_dst_eretaddr~1 .extended_lut = "off";
defparam \D_ctrl_implicit_dst_eretaddr~1 .lut_mask = 64'hFFFFFFFFBBF3FFFF;
defparam \D_ctrl_implicit_dst_eretaddr~1 .shared_arith = "off";

dffeas \W_alu_result[4] (
	.clk(clk_clk),
	.d(\E_alu_result[4]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_4),
	.prn(vcc));
defparam \W_alu_result[4] .is_wysiwyg = "true";
defparam \W_alu_result[4] .power_up = "low";

dffeas \W_alu_result[11] (
	.clk(clk_clk),
	.d(\E_alu_result[11]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_11),
	.prn(vcc));
defparam \W_alu_result[11] .is_wysiwyg = "true";
defparam \W_alu_result[11] .power_up = "low";

dffeas \W_alu_result[10] (
	.clk(clk_clk),
	.d(\E_alu_result[10]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_10),
	.prn(vcc));
defparam \W_alu_result[10] .is_wysiwyg = "true";
defparam \W_alu_result[10] .power_up = "low";

dffeas \W_alu_result[9] (
	.clk(clk_clk),
	.d(\E_alu_result[9]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_9),
	.prn(vcc));
defparam \W_alu_result[9] .is_wysiwyg = "true";
defparam \W_alu_result[9] .power_up = "low";

dffeas \W_alu_result[8] (
	.clk(clk_clk),
	.d(\E_alu_result[8]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_8),
	.prn(vcc));
defparam \W_alu_result[8] .is_wysiwyg = "true";
defparam \W_alu_result[8] .power_up = "low";

dffeas \W_alu_result[7] (
	.clk(clk_clk),
	.d(\E_alu_result[7]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_7),
	.prn(vcc));
defparam \W_alu_result[7] .is_wysiwyg = "true";
defparam \W_alu_result[7] .power_up = "low";

dffeas \W_alu_result[6] (
	.clk(clk_clk),
	.d(\E_alu_result[6]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_6),
	.prn(vcc));
defparam \W_alu_result[6] .is_wysiwyg = "true";
defparam \W_alu_result[6] .power_up = "low";

dffeas \W_alu_result[5] (
	.clk(clk_clk),
	.d(\E_alu_result[5]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_5),
	.prn(vcc));
defparam \W_alu_result[5] .is_wysiwyg = "true";
defparam \W_alu_result[5] .power_up = "low";

dffeas \W_alu_result[12] (
	.clk(clk_clk),
	.d(\E_alu_result[12]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_12),
	.prn(vcc));
defparam \W_alu_result[12] .is_wysiwyg = "true";
defparam \W_alu_result[12] .power_up = "low";

dffeas \W_alu_result[13] (
	.clk(clk_clk),
	.d(\E_alu_result[13]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_13),
	.prn(vcc));
defparam \W_alu_result[13] .is_wysiwyg = "true";
defparam \W_alu_result[13] .power_up = "low";

dffeas \W_alu_result[14] (
	.clk(clk_clk),
	.d(\E_alu_result[14]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_14),
	.prn(vcc));
defparam \W_alu_result[14] .is_wysiwyg = "true";
defparam \W_alu_result[14] .power_up = "low";

dffeas \W_alu_result[15] (
	.clk(clk_clk),
	.d(\E_alu_result[15]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_15),
	.prn(vcc));
defparam \W_alu_result[15] .is_wysiwyg = "true";
defparam \W_alu_result[15] .power_up = "low";

dffeas \W_alu_result[16] (
	.clk(clk_clk),
	.d(\E_alu_result[16]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_16),
	.prn(vcc));
defparam \W_alu_result[16] .is_wysiwyg = "true";
defparam \W_alu_result[16] .power_up = "low";

dffeas \W_alu_result[3] (
	.clk(clk_clk),
	.d(\E_alu_result[3]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_3),
	.prn(vcc));
defparam \W_alu_result[3] .is_wysiwyg = "true";
defparam \W_alu_result[3] .power_up = "low";

dffeas \W_alu_result[2] (
	.clk(clk_clk),
	.d(\E_alu_result[2]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(W_alu_result_2),
	.prn(vcc));
defparam \W_alu_result[2] .is_wysiwyg = "true";
defparam \W_alu_result[2] .power_up = "low";

dffeas \F_pc[9] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[9]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_9),
	.prn(vcc));
defparam \F_pc[9] .is_wysiwyg = "true";
defparam \F_pc[9] .power_up = "low";

dffeas \F_pc[10] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[10]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_10),
	.prn(vcc));
defparam \F_pc[10] .is_wysiwyg = "true";
defparam \F_pc[10] .power_up = "low";

dffeas \F_pc[11] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[11]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_11),
	.prn(vcc));
defparam \F_pc[11] .is_wysiwyg = "true";
defparam \F_pc[11] .power_up = "low";

dffeas \F_pc[12] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[12]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_12),
	.prn(vcc));
defparam \F_pc[12] .is_wysiwyg = "true";
defparam \F_pc[12] .power_up = "low";

dffeas \F_pc[14] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[14]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_14),
	.prn(vcc));
defparam \F_pc[14] .is_wysiwyg = "true";
defparam \F_pc[14] .power_up = "low";

dffeas \F_pc[2] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[2]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_2),
	.prn(vcc));
defparam \F_pc[2] .is_wysiwyg = "true";
defparam \F_pc[2] .power_up = "low";

dffeas \F_pc[8] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[8]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_8),
	.prn(vcc));
defparam \F_pc[8] .is_wysiwyg = "true";
defparam \F_pc[8] .power_up = "low";

dffeas \F_pc[7] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[7]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_7),
	.prn(vcc));
defparam \F_pc[7] .is_wysiwyg = "true";
defparam \F_pc[7] .power_up = "low";

dffeas \F_pc[6] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[6]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_6),
	.prn(vcc));
defparam \F_pc[6] .is_wysiwyg = "true";
defparam \F_pc[6] .power_up = "low";

dffeas \F_pc[5] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[5]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_5),
	.prn(vcc));
defparam \F_pc[5] .is_wysiwyg = "true";
defparam \F_pc[5] .power_up = "low";

dffeas \F_pc[4] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[4]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_4),
	.prn(vcc));
defparam \F_pc[4] .is_wysiwyg = "true";
defparam \F_pc[4] .power_up = "low";

dffeas \F_pc[3] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_ctrl_exception~q ),
	.ena(\W_valid~q ),
	.q(F_pc_3),
	.prn(vcc));
defparam \F_pc[3] .is_wysiwyg = "true";
defparam \F_pc[3] .power_up = "low";

dffeas \F_pc[1] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[1]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_1),
	.prn(vcc));
defparam \F_pc[1] .is_wysiwyg = "true";
defparam \F_pc[1] .power_up = "low";

dffeas \F_pc[0] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[0]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_ctrl_exception~q ),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_0),
	.prn(vcc));
defparam \F_pc[0] .is_wysiwyg = "true";
defparam \F_pc[0] .power_up = "low";

dffeas \d_writedata[22] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(vcc),
	.q(d_writedata_22),
	.prn(vcc));
defparam \d_writedata[22] .is_wysiwyg = "true";
defparam \d_writedata[22] .power_up = "low";

dffeas \d_writedata[23] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(vcc),
	.q(d_writedata_23),
	.prn(vcc));
defparam \d_writedata[23] .is_wysiwyg = "true";
defparam \d_writedata[23] .power_up = "low";

dffeas \d_writedata[11] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_11),
	.prn(vcc));
defparam \d_writedata[11] .is_wysiwyg = "true";
defparam \d_writedata[11] .power_up = "low";

dffeas \d_writedata[12] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_12),
	.prn(vcc));
defparam \d_writedata[12] .is_wysiwyg = "true";
defparam \d_writedata[12] .power_up = "low";

dffeas \d_writedata[13] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_13),
	.prn(vcc));
defparam \d_writedata[13] .is_wysiwyg = "true";
defparam \d_writedata[13] .power_up = "low";

dffeas \d_writedata[14] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_14),
	.prn(vcc));
defparam \d_writedata[14] .is_wysiwyg = "true";
defparam \d_writedata[14] .power_up = "low";

dffeas \d_writedata[15] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_15),
	.prn(vcc));
defparam \d_writedata[15] .is_wysiwyg = "true";
defparam \d_writedata[15] .power_up = "low";

dffeas \d_writedata[16] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(vcc),
	.q(d_writedata_16),
	.prn(vcc));
defparam \d_writedata[16] .is_wysiwyg = "true";
defparam \d_writedata[16] .power_up = "low";

dffeas \d_writedata[8] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_8),
	.prn(vcc));
defparam \d_writedata[8] .is_wysiwyg = "true";
defparam \d_writedata[8] .power_up = "low";

dffeas \d_writedata[10] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_10),
	.prn(vcc));
defparam \d_writedata[10] .is_wysiwyg = "true";
defparam \d_writedata[10] .power_up = "low";

dffeas \d_writedata[17] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(vcc),
	.q(d_writedata_17),
	.prn(vcc));
defparam \d_writedata[17] .is_wysiwyg = "true";
defparam \d_writedata[17] .power_up = "low";

dffeas \d_writedata[9] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_9),
	.prn(vcc));
defparam \d_writedata[9] .is_wysiwyg = "true";
defparam \d_writedata[9] .power_up = "low";

dffeas \d_writedata[18] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(vcc),
	.q(d_writedata_18),
	.prn(vcc));
defparam \d_writedata[18] .is_wysiwyg = "true";
defparam \d_writedata[18] .power_up = "low";

dffeas \d_writedata[19] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(vcc),
	.q(d_writedata_19),
	.prn(vcc));
defparam \d_writedata[19] .is_wysiwyg = "true";
defparam \d_writedata[19] .power_up = "low";

dffeas \d_writedata[20] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(vcc),
	.q(d_writedata_20),
	.prn(vcc));
defparam \d_writedata[20] .is_wysiwyg = "true";
defparam \d_writedata[20] .power_up = "low";

dffeas \d_writedata[21] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_st_data[23]~0_combout ),
	.ena(vcc),
	.q(d_writedata_21),
	.prn(vcc));
defparam \d_writedata[21] .is_wysiwyg = "true";
defparam \d_writedata[21] .power_up = "low";

dffeas \d_writedata[0] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_0),
	.prn(vcc));
defparam \d_writedata[0] .is_wysiwyg = "true";
defparam \d_writedata[0] .power_up = "low";

dffeas d_write(
	.clk(clk_clk),
	.d(\E_st_stall~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_write1),
	.prn(vcc));
defparam d_write.is_wysiwyg = "true";
defparam d_write.power_up = "low";

dffeas \d_writedata[1] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_1),
	.prn(vcc));
defparam \d_writedata[1] .is_wysiwyg = "true";
defparam \d_writedata[1] .power_up = "low";

dffeas \d_writedata[2] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_2),
	.prn(vcc));
defparam \d_writedata[2] .is_wysiwyg = "true";
defparam \d_writedata[2] .power_up = "low";

dffeas \d_writedata[3] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_3),
	.prn(vcc));
defparam \d_writedata[3] .is_wysiwyg = "true";
defparam \d_writedata[3] .power_up = "low";

dffeas \d_writedata[4] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_4),
	.prn(vcc));
defparam \d_writedata[4] .is_wysiwyg = "true";
defparam \d_writedata[4] .power_up = "low";

dffeas \d_writedata[5] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_5),
	.prn(vcc));
defparam \d_writedata[5] .is_wysiwyg = "true";
defparam \d_writedata[5] .power_up = "low";

dffeas d_read(
	.clk(clk_clk),
	.d(\d_read_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_read1),
	.prn(vcc));
defparam d_read.is_wysiwyg = "true";
defparam d_read.power_up = "low";

dffeas i_read(
	.clk(clk_clk),
	.d(\i_read_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(i_read1),
	.prn(vcc));
defparam i_read.is_wysiwyg = "true";
defparam i_read.power_up = "low";

dffeas \F_pc[13] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[13]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_13),
	.prn(vcc));
defparam \F_pc[13] .is_wysiwyg = "true";
defparam \F_pc[13] .power_up = "low";

dffeas hbreak_enabled(
	.clk(clk_clk),
	.d(\hbreak_enabled~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(hbreak_enabled1),
	.prn(vcc));
defparam hbreak_enabled.is_wysiwyg = "true";
defparam hbreak_enabled.power_up = "low";

dffeas \d_byteenable[0] (
	.clk(clk_clk),
	.d(\E_mem_byte_en~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_0),
	.prn(vcc));
defparam \d_byteenable[0] .is_wysiwyg = "true";
defparam \d_byteenable[0] .power_up = "low";

dffeas \d_byteenable[2] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_2),
	.prn(vcc));
defparam \d_byteenable[2] .is_wysiwyg = "true";
defparam \d_byteenable[2] .power_up = "low";

dffeas \d_writedata[24] (
	.clk(clk_clk),
	.d(\E_st_data[24]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_24),
	.prn(vcc));
defparam \d_writedata[24] .is_wysiwyg = "true";
defparam \d_writedata[24] .power_up = "low";

dffeas \d_byteenable[3] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[3]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_3),
	.prn(vcc));
defparam \d_byteenable[3] .is_wysiwyg = "true";
defparam \d_byteenable[3] .power_up = "low";

dffeas \d_writedata[25] (
	.clk(clk_clk),
	.d(\E_st_data[25]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_25),
	.prn(vcc));
defparam \d_writedata[25] .is_wysiwyg = "true";
defparam \d_writedata[25] .power_up = "low";

dffeas \d_writedata[26] (
	.clk(clk_clk),
	.d(\E_st_data[26]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_26),
	.prn(vcc));
defparam \d_writedata[26] .is_wysiwyg = "true";
defparam \d_writedata[26] .power_up = "low";

dffeas \d_byteenable[1] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[1]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_1),
	.prn(vcc));
defparam \d_byteenable[1] .is_wysiwyg = "true";
defparam \d_byteenable[1] .power_up = "low";

dffeas \d_writedata[6] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_6),
	.prn(vcc));
defparam \d_writedata[6] .is_wysiwyg = "true";
defparam \d_writedata[6] .power_up = "low";

dffeas \d_writedata[7] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_7),
	.prn(vcc));
defparam \d_writedata[7] .is_wysiwyg = "true";
defparam \d_writedata[7] .power_up = "low";

dffeas \d_writedata[27] (
	.clk(clk_clk),
	.d(\E_st_data[27]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_27),
	.prn(vcc));
defparam \d_writedata[27] .is_wysiwyg = "true";
defparam \d_writedata[27] .power_up = "low";

dffeas \d_writedata[28] (
	.clk(clk_clk),
	.d(\E_st_data[28]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_28),
	.prn(vcc));
defparam \d_writedata[28] .is_wysiwyg = "true";
defparam \d_writedata[28] .power_up = "low";

dffeas \d_writedata[29] (
	.clk(clk_clk),
	.d(\E_st_data[29]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_29),
	.prn(vcc));
defparam \d_writedata[29] .is_wysiwyg = "true";
defparam \d_writedata[29] .power_up = "low";

dffeas \d_writedata[30] (
	.clk(clk_clk),
	.d(\E_st_data[30]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_30),
	.prn(vcc));
defparam \d_writedata[30] .is_wysiwyg = "true";
defparam \d_writedata[30] .power_up = "low";

dffeas \d_writedata[31] (
	.clk(clk_clk),
	.d(\E_st_data[31]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_31),
	.prn(vcc));
defparam \d_writedata[31] .is_wysiwyg = "true";
defparam \d_writedata[31] .power_up = "low";

cyclonev_lcell_comb \F_valid~0 (
	.dataa(!i_read1),
	.datab(!src1_valid1),
	.datac(!src1_valid2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_valid~0 .extended_lut = "off";
defparam \F_valid~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \F_valid~0 .shared_arith = "off";

dffeas D_valid(
	.clk(clk_clk),
	.d(\F_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\D_valid~q ),
	.prn(vcc));
defparam D_valid.is_wysiwyg = "true";
defparam D_valid.power_up = "low";

dffeas R_valid(
	.clk(clk_clk),
	.d(\D_valid~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_valid~q ),
	.prn(vcc));
defparam R_valid.is_wysiwyg = "true";
defparam R_valid.power_up = "low";

dffeas E_new_inst(
	.clk(clk_clk),
	.d(\R_valid~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_new_inst~q ),
	.prn(vcc));
defparam E_new_inst.is_wysiwyg = "true";
defparam E_new_inst.power_up = "low";

dffeas \D_iw[0] (
	.clk(clk_clk),
	.d(src_data_01),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[0]~q ),
	.prn(vcc));
defparam \D_iw[0] .is_wysiwyg = "true";
defparam \D_iw[0] .power_up = "low";

cyclonev_lcell_comb \F_iw[1]~4 (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!av_readdata_pre_1),
	.datad(!q_a_1),
	.datae(!\hbreak_req~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[1]~4 .extended_lut = "off";
defparam \F_iw[1]~4 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \F_iw[1]~4 .shared_arith = "off";

dffeas \D_iw[1] (
	.clk(clk_clk),
	.d(\F_iw[1]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[1]~q ),
	.prn(vcc));
defparam \D_iw[1] .is_wysiwyg = "true";
defparam \D_iw[1] .power_up = "low";

cyclonev_lcell_comb \F_iw[4]~6 (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!av_readdata_pre_4),
	.datad(!q_a_4),
	.datae(!\hbreak_req~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[4]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[4]~6 .extended_lut = "off";
defparam \F_iw[4]~6 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \F_iw[4]~6 .shared_arith = "off";

dffeas \D_iw[4] (
	.clk(clk_clk),
	.d(\F_iw[4]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[4]~q ),
	.prn(vcc));
defparam \D_iw[4] .is_wysiwyg = "true";
defparam \D_iw[4] .power_up = "low";

cyclonev_lcell_comb \F_iw[3]~5 (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!av_readdata_pre_3),
	.datad(!q_a_3),
	.datae(!\hbreak_req~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[3]~5 .extended_lut = "off";
defparam \F_iw[3]~5 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \F_iw[3]~5 .shared_arith = "off";

dffeas \D_iw[3] (
	.clk(clk_clk),
	.d(\F_iw[3]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[3]~q ),
	.prn(vcc));
defparam \D_iw[3] .is_wysiwyg = "true";
defparam \D_iw[3] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_st~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[4]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_st~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_st~0 .extended_lut = "off";
defparam \D_ctrl_st~0 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \D_ctrl_st~0 .shared_arith = "off";

dffeas \D_iw[2] (
	.clk(clk_clk),
	.d(src_data_2),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[2]~q ),
	.prn(vcc));
defparam \D_iw[2] .is_wysiwyg = "true";
defparam \D_iw[2] .power_up = "low";

dffeas R_ctrl_st(
	.clk(clk_clk),
	.d(\D_ctrl_st~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!\D_iw[2]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_st~q ),
	.prn(vcc));
defparam R_ctrl_st.is_wysiwyg = "true";
defparam R_ctrl_st.power_up = "low";

cyclonev_lcell_comb \d_write_nxt~0 (
	.dataa(!\E_new_inst~q ),
	.datab(!\R_ctrl_st~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_write_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_write_nxt~0 .extended_lut = "off";
defparam \d_write_nxt~0 .lut_mask = 64'h7777777777777777;
defparam \d_write_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_ld~0 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_ld~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_ld~0 .extended_lut = "off";
defparam \D_ctrl_ld~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \D_ctrl_ld~0 .shared_arith = "off";

dffeas R_ctrl_ld(
	.clk(clk_clk),
	.d(\D_ctrl_ld~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_ld~q ),
	.prn(vcc));
defparam R_ctrl_ld.is_wysiwyg = "true";
defparam R_ctrl_ld.power_up = "low";

dffeas av_ld_waiting_for_data(
	.clk(clk_clk),
	.d(\av_ld_waiting_for_data_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_waiting_for_data~q ),
	.prn(vcc));
defparam av_ld_waiting_for_data.is_wysiwyg = "true";
defparam av_ld_waiting_for_data.power_up = "low";

cyclonev_lcell_comb \av_ld_waiting_for_data_nxt~0 (
	.dataa(!d_read1),
	.datab(!\E_new_inst~q ),
	.datac(!src0_valid),
	.datad(!WideOr1),
	.datae(!\R_ctrl_ld~q ),
	.dataf(!\av_ld_waiting_for_data~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_waiting_for_data_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_waiting_for_data_nxt~0 .extended_lut = "off";
defparam \av_ld_waiting_for_data_nxt~0 .lut_mask = 64'hBBFFFFFFF3FFFFFF;
defparam \av_ld_waiting_for_data_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_mem32~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[2]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_mem32~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_mem32~0 .extended_lut = "off";
defparam \D_ctrl_mem32~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \D_ctrl_mem32~0 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_aligning_data_nxt~1 (
	.dataa(!d_read1),
	.datab(!src0_valid),
	.datac(!WideOr1),
	.datad(!\av_ld_aligning_data~q ),
	.datae(!\D_ctrl_mem32~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_aligning_data_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_aligning_data_nxt~1 .extended_lut = "off";
defparam \av_ld_aligning_data_nxt~1 .lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam \av_ld_aligning_data_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_aligning_data_nxt~2 (
	.dataa(!\av_ld_aligning_data_nxt~0_combout ),
	.datab(!\av_ld_aligning_data_nxt~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_aligning_data_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_aligning_data_nxt~2 .extended_lut = "off";
defparam \av_ld_aligning_data_nxt~2 .lut_mask = 64'h7777777777777777;
defparam \av_ld_aligning_data_nxt~2 .shared_arith = "off";

dffeas av_ld_aligning_data(
	.clk(clk_clk),
	.d(\av_ld_aligning_data_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_aligning_data~q ),
	.prn(vcc));
defparam av_ld_aligning_data.is_wysiwyg = "true";
defparam av_ld_aligning_data.power_up = "low";

cyclonev_lcell_comb \av_ld_align_cycle_nxt[0]~1 (
	.dataa(!d_read1),
	.datab(!src0_valid),
	.datac(!WideOr1),
	.datad(!\av_ld_align_cycle[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_align_cycle_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_align_cycle_nxt[0]~1 .extended_lut = "off";
defparam \av_ld_align_cycle_nxt[0]~1 .lut_mask = 64'hFFEFFFEFFFEFFFEF;
defparam \av_ld_align_cycle_nxt[0]~1 .shared_arith = "off";

dffeas \av_ld_align_cycle[0] (
	.clk(clk_clk),
	.d(\av_ld_align_cycle_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_align_cycle[0]~q ),
	.prn(vcc));
defparam \av_ld_align_cycle[0] .is_wysiwyg = "true";
defparam \av_ld_align_cycle[0] .power_up = "low";

cyclonev_lcell_comb \av_ld_align_cycle_nxt[1]~0 (
	.dataa(!d_read1),
	.datab(!src0_valid),
	.datac(!WideOr1),
	.datad(!\av_ld_align_cycle[1]~q ),
	.datae(!\av_ld_align_cycle[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_align_cycle_nxt[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_align_cycle_nxt[1]~0 .extended_lut = "off";
defparam \av_ld_align_cycle_nxt[1]~0 .lut_mask = 64'hEFFFFFEFEFFFFFEF;
defparam \av_ld_align_cycle_nxt[1]~0 .shared_arith = "off";

dffeas \av_ld_align_cycle[1] (
	.clk(clk_clk),
	.d(\av_ld_align_cycle_nxt[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_align_cycle[1]~q ),
	.prn(vcc));
defparam \av_ld_align_cycle[1] .is_wysiwyg = "true";
defparam \av_ld_align_cycle[1] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_mem16~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_mem16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_mem16~0 .extended_lut = "off";
defparam \D_ctrl_mem16~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_ctrl_mem16~0 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_aligning_data_nxt~0 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\av_ld_aligning_data~q ),
	.datac(!\av_ld_align_cycle[1]~q ),
	.datad(!\av_ld_align_cycle[0]~q ),
	.datae(!\D_ctrl_mem16~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_aligning_data_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_aligning_data_nxt~0 .extended_lut = "off";
defparam \av_ld_aligning_data_nxt~0 .lut_mask = 64'hFBF7F7FBFBF7F7FB;
defparam \av_ld_aligning_data_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \E_ld_stall~0 (
	.dataa(!\R_ctrl_ld~q ),
	.datab(!\E_valid_from_R~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ld_stall~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ld_stall~0 .extended_lut = "off";
defparam \E_ld_stall~0 .lut_mask = 64'h7777777777777777;
defparam \E_ld_stall~0 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[5]~7 (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!av_readdata_pre_5),
	.datad(!q_a_5),
	.datae(!\hbreak_req~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[5]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[5]~7 .extended_lut = "off";
defparam \F_iw[5]~7 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \F_iw[5]~7 .shared_arith = "off";

dffeas \D_iw[5] (
	.clk(clk_clk),
	.d(\F_iw[5]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[5]~q ),
	.prn(vcc));
defparam \D_iw[5] .is_wysiwyg = "true";
defparam \D_iw[5] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_b_is_dst~0 (
	.dataa(!\D_iw[3]~q ),
	.datab(!\D_iw[2]~q ),
	.datac(!\D_iw[1]~q ),
	.datad(!\D_iw[0]~q ),
	.datae(!\D_iw[5]~q ),
	.dataf(!\D_iw[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_b_is_dst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_b_is_dst~0 .extended_lut = "off";
defparam \D_ctrl_b_is_dst~0 .lut_mask = 64'hFFFF9669FFFF6996;
defparam \D_ctrl_b_is_dst~0 .shared_arith = "off";

cyclonev_lcell_comb \R_ctrl_br_nxt~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[5]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_ctrl_br_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_ctrl_br_nxt~0 .extended_lut = "off";
defparam \R_ctrl_br_nxt~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \R_ctrl_br_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \R_ctrl_br_nxt~1 (
	.dataa(!\D_iw[1]~q ),
	.datab(!\D_iw[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_ctrl_br_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_ctrl_br_nxt~1 .extended_lut = "off";
defparam \R_ctrl_br_nxt~1 .lut_mask = 64'h7777777777777777;
defparam \R_ctrl_br_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \R_ctrl_br_nxt~2 (
	.dataa(!\R_ctrl_br_nxt~0_combout ),
	.datab(!\R_ctrl_br_nxt~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_ctrl_br_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_ctrl_br_nxt~2 .extended_lut = "off";
defparam \R_ctrl_br_nxt~2 .lut_mask = 64'h7777777777777777;
defparam \R_ctrl_br_nxt~2 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[13]~1 (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!av_readdata_pre_13),
	.datad(!q_a_13),
	.datae(!\hbreak_req~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[13]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[13]~1 .extended_lut = "off";
defparam \F_iw[13]~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \F_iw[13]~1 .shared_arith = "off";

dffeas \D_iw[13] (
	.clk(clk_clk),
	.d(\F_iw[13]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[13]~q ),
	.prn(vcc));
defparam \D_iw[13] .is_wysiwyg = "true";
defparam \D_iw[13] .power_up = "low";

dffeas \D_iw[12] (
	.clk(clk_clk),
	.d(src_data_12),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[12]~q ),
	.prn(vcc));
defparam \D_iw[12] .is_wysiwyg = "true";
defparam \D_iw[12] .power_up = "low";

cyclonev_lcell_comb \F_iw[15]~2 (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!av_readdata_pre_15),
	.datad(!q_a_15),
	.datae(!\hbreak_req~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[15]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[15]~2 .extended_lut = "off";
defparam \F_iw[15]~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \F_iw[15]~2 .shared_arith = "off";

dffeas \D_iw[15] (
	.clk(clk_clk),
	.d(\F_iw[15]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[15]~q ),
	.prn(vcc));
defparam \D_iw[15] .is_wysiwyg = "true";
defparam \D_iw[15] .power_up = "low";

cyclonev_lcell_comb \F_iw[11]~0 (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!av_readdata_pre_11),
	.datad(!q_a_11),
	.datae(!\hbreak_req~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[11]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[11]~0 .extended_lut = "off";
defparam \F_iw[11]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \F_iw[11]~0 .shared_arith = "off";

dffeas \D_iw[11] (
	.clk(clk_clk),
	.d(\F_iw[11]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[11]~q ),
	.prn(vcc));
defparam \D_iw[11] .is_wysiwyg = "true";
defparam \D_iw[11] .power_up = "low";

dffeas \D_iw[14] (
	.clk(clk_clk),
	.d(src_data_14),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[14]~q ),
	.prn(vcc));
defparam \D_iw[14] .is_wysiwyg = "true";
defparam \D_iw[14] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hFBFFFFFFFFFFFFFF;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \R_src2_use_imm~1 (
	.dataa(!\D_iw[13]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[15]~q ),
	.datad(!\D_iw[11]~q ),
	.datae(!\D_iw[14]~q ),
	.dataf(!\Equal0~0_combout ),
	.datag(!\D_iw[16]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_use_imm~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_use_imm~1 .extended_lut = "on";
defparam \R_src2_use_imm~1 .lut_mask = 64'hDFFFFDFFDFFFFDFF;
defparam \R_src2_use_imm~1 .shared_arith = "off";

cyclonev_lcell_comb \R_src2_use_imm~5 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_use_imm~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_use_imm~5 .extended_lut = "off";
defparam \R_src2_use_imm~5 .lut_mask = 64'hFFEFFFFFFFEFFFFF;
defparam \R_src2_use_imm~5 .shared_arith = "off";

cyclonev_lcell_comb \R_src2_use_imm~0 (
	.dataa(!\R_valid~q ),
	.datab(!\D_ctrl_b_is_dst~0_combout ),
	.datac(!\R_ctrl_br_nxt~2_combout ),
	.datad(!\R_src2_use_imm~1_combout ),
	.datae(!\R_src2_use_imm~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_use_imm~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_use_imm~0 .extended_lut = "off";
defparam \R_src2_use_imm~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \R_src2_use_imm~0 .shared_arith = "off";

dffeas R_src2_use_imm(
	.clk(clk_clk),
	.d(\R_src2_use_imm~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_src2_use_imm~q ),
	.prn(vcc));
defparam R_src2_use_imm.is_wysiwyg = "true";
defparam R_src2_use_imm.power_up = "low";

cyclonev_lcell_comb \D_ctrl_src_imm5_shift_rot~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[16]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_src_imm5_shift_rot~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_src_imm5_shift_rot~0 .extended_lut = "off";
defparam \D_ctrl_src_imm5_shift_rot~0 .lut_mask = 64'hBBF3BBF3BBF3BBF3;
defparam \D_ctrl_src_imm5_shift_rot~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_src_imm5_shift_rot~1 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\Equal0~0_combout ),
	.datad(!\D_ctrl_src_imm5_shift_rot~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_src_imm5_shift_rot~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_src_imm5_shift_rot~1 .extended_lut = "off";
defparam \D_ctrl_src_imm5_shift_rot~1 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \D_ctrl_src_imm5_shift_rot~1 .shared_arith = "off";

dffeas R_ctrl_src_imm5_shift_rot(
	.clk(clk_clk),
	.d(\D_ctrl_src_imm5_shift_rot~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_src_imm5_shift_rot~q ),
	.prn(vcc));
defparam R_ctrl_src_imm5_shift_rot.is_wysiwyg = "true";
defparam R_ctrl_src_imm5_shift_rot.power_up = "low";

cyclonev_lcell_comb \R_src2_lo~0 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\R_ctrl_src_imm5_shift_rot~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_lo~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_lo~0 .extended_lut = "off";
defparam \R_src2_lo~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \R_src2_lo~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_hi_imm16~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[4]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[2]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_hi_imm16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_hi_imm16~0 .extended_lut = "off";
defparam \D_ctrl_hi_imm16~0 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \D_ctrl_hi_imm16~0 .shared_arith = "off";

dffeas R_ctrl_hi_imm16(
	.clk(clk_clk),
	.d(\D_ctrl_hi_imm16~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_hi_imm16~q ),
	.prn(vcc));
defparam R_ctrl_hi_imm16.is_wysiwyg = "true";
defparam R_ctrl_hi_imm16.power_up = "low";

cyclonev_lcell_comb \Equal62~7 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~7 .extended_lut = "off";
defparam \Equal62~7 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \Equal62~7 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~8 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~8 .extended_lut = "off";
defparam \Equal62~8 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \Equal62~8 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_implicit_dst_eretaddr~5 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_implicit_dst_eretaddr~5 .extended_lut = "off";
defparam \D_ctrl_implicit_dst_eretaddr~5 .lut_mask = 64'hD77D7DD77DD7D77D;
defparam \D_ctrl_implicit_dst_eretaddr~5 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_implicit_dst_eretaddr~4 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_implicit_dst_eretaddr~4 .extended_lut = "off";
defparam \D_ctrl_implicit_dst_eretaddr~4 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \D_ctrl_implicit_dst_eretaddr~4 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_implicit_dst_eretaddr~3 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_implicit_dst_eretaddr~3 .extended_lut = "off";
defparam \D_ctrl_implicit_dst_eretaddr~3 .lut_mask = 64'hFF69FF96FFFFFFFF;
defparam \D_ctrl_implicit_dst_eretaddr~3 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_implicit_dst_eretaddr~0 (
	.dataa(!\Equal62~7_combout ),
	.datab(!\Equal62~8_combout ),
	.datac(!\D_ctrl_implicit_dst_eretaddr~5_combout ),
	.datad(!\D_ctrl_implicit_dst_eretaddr~4_combout ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_implicit_dst_eretaddr~0 .extended_lut = "off";
defparam \D_ctrl_implicit_dst_eretaddr~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \D_ctrl_implicit_dst_eretaddr~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~10 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~10 .extended_lut = "off";
defparam \Equal0~10 .lut_mask = 64'hFFFFFBFFFFFFFFFF;
defparam \Equal0~10 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_exception~6 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_exception~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_exception~6 .extended_lut = "off";
defparam \D_ctrl_exception~6 .lut_mask = 64'h7FFFFF7FFFFFFFFF;
defparam \D_ctrl_exception~6 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_exception~5 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_exception~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_exception~5 .extended_lut = "off";
defparam \D_ctrl_exception~5 .lut_mask = 64'hFFBFFFFFFFFFFFBF;
defparam \D_ctrl_exception~5 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_exception~4 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_exception~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_exception~4 .extended_lut = "off";
defparam \D_ctrl_exception~4 .lut_mask = 64'h6996966996696996;
defparam \D_ctrl_exception~4 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_exception~1 (
	.dataa(!\Equal0~10_combout ),
	.datab(!\D_ctrl_exception~6_combout ),
	.datac(!\D_ctrl_exception~5_combout ),
	.datad(!\D_ctrl_exception~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_exception~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_exception~1 .extended_lut = "off";
defparam \D_ctrl_exception~1 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \D_ctrl_exception~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~9 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~9 .extended_lut = "off";
defparam \Equal62~9 .lut_mask = 64'hFFEFFFFFFFFFFFFF;
defparam \Equal62~9 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~10 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~10 .extended_lut = "off";
defparam \Equal62~10 .lut_mask = 64'hFFDFFFFFFFFFFFFF;
defparam \Equal62~10 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~11 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~11 .extended_lut = "off";
defparam \Equal62~11 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \Equal62~11 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~13 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~13 .extended_lut = "off";
defparam \Equal62~13 .lut_mask = 64'hFFFFFFFFFFFFFFDF;
defparam \Equal62~13 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~14 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~14 .extended_lut = "off";
defparam \Equal62~14 .lut_mask = 64'hFFFFFFFFFFFFDFFF;
defparam \Equal62~14 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_force_src2_zero~0 (
	.dataa(!\Equal62~9_combout ),
	.datab(!\Equal62~10_combout ),
	.datac(!\Equal62~11_combout ),
	.datad(!\Equal62~13_combout ),
	.datae(!\Equal62~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_force_src2_zero~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_force_src2_zero~0 .extended_lut = "off";
defparam \D_ctrl_force_src2_zero~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \D_ctrl_force_src2_zero~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~7 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~7 .extended_lut = "off";
defparam \Equal0~7 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal0~7 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~8 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~8 .extended_lut = "off";
defparam \Equal0~8 .lut_mask = 64'hFFFFFFFFFFFFFFFB;
defparam \Equal0~8 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_retaddr~2 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_retaddr~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_retaddr~2 .extended_lut = "off";
defparam \D_ctrl_retaddr~2 .lut_mask = 64'hFFFF6FFFFFFF6FFF;
defparam \D_ctrl_retaddr~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_retaddr~0 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal0~7_combout ),
	.datac(!\Equal0~8_combout ),
	.datad(!\D_ctrl_retaddr~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_retaddr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_retaddr~0 .extended_lut = "off";
defparam \D_ctrl_retaddr~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \D_ctrl_retaddr~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~11 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~11 .extended_lut = "off";
defparam \Equal0~11 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \Equal0~11 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~15 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~15 .extended_lut = "off";
defparam \Equal62~15 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \Equal62~15 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~16 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~16 .extended_lut = "off";
defparam \Equal62~16 .lut_mask = 64'hFFFFFFFFFFFFFDFF;
defparam \Equal62~16 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_force_src2_zero~1 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal0~11_combout ),
	.datac(!\Equal62~15_combout ),
	.datad(!\Equal62~16_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_force_src2_zero~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_force_src2_zero~1 .extended_lut = "off";
defparam \D_ctrl_force_src2_zero~1 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \D_ctrl_force_src2_zero~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_force_src2_zero~2 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.datac(!\D_ctrl_exception~1_combout ),
	.datad(!\D_ctrl_force_src2_zero~0_combout ),
	.datae(!\D_ctrl_retaddr~0_combout ),
	.dataf(!\D_ctrl_force_src2_zero~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_force_src2_zero~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_force_src2_zero~2 .extended_lut = "off";
defparam \D_ctrl_force_src2_zero~2 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \D_ctrl_force_src2_zero~2 .shared_arith = "off";

dffeas R_ctrl_force_src2_zero(
	.clk(clk_clk),
	.d(\D_ctrl_force_src2_zero~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_force_src2_zero~q ),
	.prn(vcc));
defparam R_ctrl_force_src2_zero.is_wysiwyg = "true";
defparam R_ctrl_force_src2_zero.power_up = "low";

dffeas \D_iw[6] (
	.clk(clk_clk),
	.d(src_data_6),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[6]~q ),
	.prn(vcc));
defparam \D_iw[6] .is_wysiwyg = "true";
defparam \D_iw[6] .power_up = "low";

cyclonev_lcell_comb \R_src2_lo[0]~5 (
	.dataa(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datab(!\R_src2_lo~0_combout ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\R_ctrl_force_src2_zero~q ),
	.datae(!\D_iw[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_lo[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_lo[0]~5 .extended_lut = "off";
defparam \R_src2_lo[0]~5 .lut_mask = 64'hF7D5FFFFF7D5FFFF;
defparam \R_src2_lo[0]~5 .shared_arith = "off";

dffeas \E_src2[0] (
	.clk(clk_clk),
	.d(\R_src2_lo[0]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[0]~q ),
	.prn(vcc));
defparam \E_src2[0] .is_wysiwyg = "true";
defparam \E_src2[0] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_cnt[0]~_wirecell (
	.dataa(!\E_shift_rot_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_cnt[0]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_cnt[0]~_wirecell .extended_lut = "off";
defparam \E_shift_rot_cnt[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \E_shift_rot_cnt[0]~_wirecell .shared_arith = "off";

dffeas \E_shift_rot_cnt[0] (
	.clk(clk_clk),
	.d(\E_src2[0]~q ),
	.asdata(\E_shift_rot_cnt[0]~_wirecell_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[0]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[0] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[0] .power_up = "low";

cyclonev_lcell_comb \Add3~3 (
	.dataa(!\E_shift_rot_cnt[1]~q ),
	.datab(!\E_shift_rot_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add3~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~3 .extended_lut = "off";
defparam \Add3~3 .lut_mask = 64'h6666666666666666;
defparam \Add3~3 .shared_arith = "off";

dffeas \D_iw[7] (
	.clk(clk_clk),
	.d(src_data_7),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[7]~q ),
	.prn(vcc));
defparam \D_iw[7] .is_wysiwyg = "true";
defparam \D_iw[7] .power_up = "low";

cyclonev_lcell_comb \R_src2_lo[1]~4 (
	.dataa(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datab(!\R_src2_lo~0_combout ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\R_ctrl_force_src2_zero~q ),
	.datae(!\D_iw[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_lo[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_lo[1]~4 .extended_lut = "off";
defparam \R_src2_lo[1]~4 .lut_mask = 64'hF7D5FFFFF7D5FFFF;
defparam \R_src2_lo[1]~4 .shared_arith = "off";

dffeas \E_src2[1] (
	.clk(clk_clk),
	.d(\R_src2_lo[1]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[1]~q ),
	.prn(vcc));
defparam \E_src2[1] .is_wysiwyg = "true";
defparam \E_src2[1] .power_up = "low";

dffeas \E_shift_rot_cnt[1] (
	.clk(clk_clk),
	.d(\Add3~3_combout ),
	.asdata(\E_src2[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[1]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[1] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[1] .power_up = "low";

cyclonev_lcell_comb \Add3~2 (
	.dataa(!\E_shift_rot_cnt[2]~q ),
	.datab(!\E_shift_rot_cnt[1]~q ),
	.datac(!\E_shift_rot_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~2 .extended_lut = "off";
defparam \Add3~2 .lut_mask = 64'h9696969696969696;
defparam \Add3~2 .shared_arith = "off";

dffeas \D_iw[8] (
	.clk(clk_clk),
	.d(src_data_8),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[8]~q ),
	.prn(vcc));
defparam \D_iw[8] .is_wysiwyg = "true";
defparam \D_iw[8] .power_up = "low";

cyclonev_lcell_comb \R_src2_lo[2]~3 (
	.dataa(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datab(!\D_iw[8]~q ),
	.datac(!\R_src2_lo~0_combout ),
	.datad(!\R_ctrl_hi_imm16~q ),
	.datae(!\R_ctrl_force_src2_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_lo[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_lo[2]~3 .extended_lut = "off";
defparam \R_src2_lo[2]~3 .lut_mask = 64'hFF7FF777FF7FF777;
defparam \R_src2_lo[2]~3 .shared_arith = "off";

dffeas \E_src2[2] (
	.clk(clk_clk),
	.d(\R_src2_lo[2]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[2]~q ),
	.prn(vcc));
defparam \E_src2[2] .is_wysiwyg = "true";
defparam \E_src2[2] .power_up = "low";

dffeas \E_shift_rot_cnt[2] (
	.clk(clk_clk),
	.d(\Add3~2_combout ),
	.asdata(\E_src2[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[2]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[2] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[2] .power_up = "low";

cyclonev_lcell_comb \Add3~1 (
	.dataa(!\E_shift_rot_cnt[3]~q ),
	.datab(!\E_shift_rot_cnt[2]~q ),
	.datac(!\E_shift_rot_cnt[1]~q ),
	.datad(!\E_shift_rot_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h6996699669966996;
defparam \Add3~1 .shared_arith = "off";

dffeas \D_iw[9] (
	.clk(clk_clk),
	.d(src_data_9),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[9]~q ),
	.prn(vcc));
defparam \D_iw[9] .is_wysiwyg = "true";
defparam \D_iw[9] .power_up = "low";

cyclonev_lcell_comb \R_src2_lo[3]~2 (
	.dataa(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datab(!\R_src2_lo~0_combout ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\R_ctrl_force_src2_zero~q ),
	.datae(!\D_iw[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_lo[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_lo[3]~2 .extended_lut = "off";
defparam \R_src2_lo[3]~2 .lut_mask = 64'hF7D5FFFFF7D5FFFF;
defparam \R_src2_lo[3]~2 .shared_arith = "off";

dffeas \E_src2[3] (
	.clk(clk_clk),
	.d(\R_src2_lo[3]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[3]~q ),
	.prn(vcc));
defparam \E_src2[3] .is_wysiwyg = "true";
defparam \E_src2[3] .power_up = "low";

dffeas \E_shift_rot_cnt[3] (
	.clk(clk_clk),
	.d(\Add3~1_combout ),
	.asdata(\E_src2[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[3]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[3] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[3] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_done~0 (
	.dataa(!\E_shift_rot_cnt[3]~q ),
	.datab(!\E_shift_rot_cnt[2]~q ),
	.datac(!\E_shift_rot_cnt[1]~q ),
	.datad(!\E_shift_rot_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_done~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_done~0 .extended_lut = "off";
defparam \E_shift_rot_done~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \E_shift_rot_done~0 .shared_arith = "off";

cyclonev_lcell_comb \Add3~0 (
	.dataa(!\E_shift_rot_cnt[4]~q ),
	.datab(!\E_shift_rot_done~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~0 .extended_lut = "off";
defparam \Add3~0 .lut_mask = 64'h6666666666666666;
defparam \Add3~0 .shared_arith = "off";

dffeas \D_iw[10] (
	.clk(clk_clk),
	.d(src_data_10),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[10]~q ),
	.prn(vcc));
defparam \D_iw[10] .is_wysiwyg = "true";
defparam \D_iw[10] .power_up = "low";

cyclonev_lcell_comb \R_src2_lo[4]~1 (
	.dataa(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datab(!\R_src2_lo~0_combout ),
	.datac(!\D_iw[10]~q ),
	.datad(!\R_ctrl_hi_imm16~q ),
	.datae(!\R_ctrl_force_src2_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_lo[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_lo[4]~1 .extended_lut = "off";
defparam \R_src2_lo[4]~1 .lut_mask = 64'hFF7FDF5FFF7FDF5F;
defparam \R_src2_lo[4]~1 .shared_arith = "off";

dffeas \E_src2[4] (
	.clk(clk_clk),
	.d(\R_src2_lo[4]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[4]~q ),
	.prn(vcc));
defparam \E_src2[4] .is_wysiwyg = "true";
defparam \E_src2[4] .power_up = "low";

dffeas \E_shift_rot_cnt[4] (
	.clk(clk_clk),
	.d(\Add3~0_combout ),
	.asdata(\E_src2[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[4]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[4] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[4] .power_up = "low";

cyclonev_lcell_comb \E_stall~0 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\E_new_inst~q ),
	.datac(!\R_ctrl_ld~q ),
	.datad(!\E_valid_from_R~q ),
	.datae(!\E_shift_rot_cnt[4]~q ),
	.dataf(!\E_shift_rot_done~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stall~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stall~0 .extended_lut = "off";
defparam \E_stall~0 .lut_mask = 64'hFFFFFFFF7FFFFFFF;
defparam \E_stall~0 .shared_arith = "off";

cyclonev_lcell_comb \E_stall~1 (
	.dataa(!\av_ld_waiting_for_data_nxt~0_combout ),
	.datab(!\av_ld_aligning_data_nxt~0_combout ),
	.datac(!\D_ctrl_mem32~0_combout ),
	.datad(!\av_ld_aligning_data_nxt~1_combout ),
	.datae(!\E_ld_stall~0_combout ),
	.dataf(!\E_stall~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stall~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stall~1 .extended_lut = "off";
defparam \E_stall~1 .lut_mask = 64'hFFFFFFFFFFFFFFEF;
defparam \E_stall~1 .shared_arith = "off";

cyclonev_lcell_comb \E_valid_from_R~0 (
	.dataa(!d_write1),
	.datab(!\d_write_nxt~0_combout ),
	.datac(!av_waitrequest2),
	.datad(!av_waitrequest),
	.datae(!\R_valid~q ),
	.dataf(!\E_stall~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_valid_from_R~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_valid_from_R~0 .extended_lut = "off";
defparam \E_valid_from_R~0 .lut_mask = 64'hFFFFFFFF7FFFFFFF;
defparam \E_valid_from_R~0 .shared_arith = "off";

dffeas E_valid_from_R(
	.clk(clk_clk),
	.d(\E_valid_from_R~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_valid_from_R~q ),
	.prn(vcc));
defparam E_valid_from_R.is_wysiwyg = "true";
defparam E_valid_from_R.power_up = "low";

cyclonev_lcell_comb \W_valid~0 (
	.dataa(!d_write1),
	.datab(!\d_write_nxt~0_combout ),
	.datac(!av_waitrequest2),
	.datad(!av_waitrequest),
	.datae(!\E_valid_from_R~q ),
	.dataf(!\E_stall~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_valid~0 .extended_lut = "off";
defparam \W_valid~0 .lut_mask = 64'hFFFEFFFFFFFFFFFF;
defparam \W_valid~0 .shared_arith = "off";

dffeas W_valid(
	.clk(clk_clk),
	.d(\W_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_valid~q ),
	.prn(vcc));
defparam W_valid.is_wysiwyg = "true";
defparam W_valid.power_up = "low";

cyclonev_lcell_comb \hbreak_pending_nxt~0 (
	.dataa(!hbreak_enabled1),
	.datab(!\hbreak_pending~q ),
	.datac(!\hbreak_req~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hbreak_pending_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hbreak_pending_nxt~0 .extended_lut = "off";
defparam \hbreak_pending_nxt~0 .lut_mask = 64'h8B8B8B8B8B8B8B8B;
defparam \hbreak_pending_nxt~0 .shared_arith = "off";

dffeas hbreak_pending(
	.clk(clk_clk),
	.d(\hbreak_pending_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\hbreak_pending~q ),
	.prn(vcc));
defparam hbreak_pending.is_wysiwyg = "true";
defparam hbreak_pending.power_up = "low";

cyclonev_lcell_comb \wait_for_one_post_bret_inst~0 (
	.dataa(!hbreak_enabled1),
	.datab(!\wait_for_one_post_bret_inst~q ),
	.datac(!\F_valid~0_combout ),
	.datad(!\the_niosLab2_nios2_gen2_0_cpu_nios2_oci|the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_for_one_post_bret_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_for_one_post_bret_inst~0 .extended_lut = "off";
defparam \wait_for_one_post_bret_inst~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \wait_for_one_post_bret_inst~0 .shared_arith = "off";

dffeas wait_for_one_post_bret_inst(
	.clk(clk_clk),
	.d(\wait_for_one_post_bret_inst~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_for_one_post_bret_inst~q ),
	.prn(vcc));
defparam wait_for_one_post_bret_inst.is_wysiwyg = "true";
defparam wait_for_one_post_bret_inst.power_up = "low";

cyclonev_lcell_comb \hbreak_req~0 (
	.dataa(!\W_valid~q ),
	.datab(!hbreak_enabled1),
	.datac(!\hbreak_pending~q ),
	.datad(!\the_niosLab2_nios2_gen2_0_cpu_nios2_oci|the_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug|jtag_break~q ),
	.datae(!\wait_for_one_post_bret_inst~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hbreak_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hbreak_req~0 .extended_lut = "off";
defparam \hbreak_req~0 .lut_mask = 64'hFFFFDFFFFFFFDFFF;
defparam \hbreak_req~0 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[16]~3 (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!av_readdata_pre_161),
	.datad(!q_a_16),
	.datae(!\hbreak_req~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[16]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[16]~3 .extended_lut = "off";
defparam \F_iw[16]~3 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \F_iw[16]~3 .shared_arith = "off";

dffeas \D_iw[16] (
	.clk(clk_clk),
	.d(\F_iw[16]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[16]~q ),
	.prn(vcc));
defparam \D_iw[16] .is_wysiwyg = "true";
defparam \D_iw[16] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_shift_rot~0 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot~0 .extended_lut = "off";
defparam \D_ctrl_shift_rot~0 .lut_mask = 64'hBFB3FFFFFFFFFFFF;
defparam \D_ctrl_shift_rot~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_shift_rot~1 (
	.dataa(gnd),
	.datab(!\D_ctrl_shift_rot~0_combout ),
	.datac(gnd),
	.datad(!\Equal0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot~1 .extended_lut = "off";
defparam \D_ctrl_shift_rot~1 .lut_mask = 64'h33FF33FF33FF33FF;
defparam \D_ctrl_shift_rot~1 .shared_arith = "off";

dffeas R_ctrl_shift_rot(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_rot~q ),
	.prn(vcc));
defparam R_ctrl_shift_rot.is_wysiwyg = "true";
defparam R_ctrl_shift_rot.power_up = "low";

cyclonev_lcell_comb \D_ctrl_shift_rot_right~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[15]~q ),
	.datad(!\D_iw[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot_right~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot_right~0 .extended_lut = "off";
defparam \D_ctrl_shift_rot_right~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \D_ctrl_shift_rot_right~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_shift_rot_right~1 (
	.dataa(!\D_iw[13]~q ),
	.datab(!\D_iw[14]~q ),
	.datac(!\Equal0~0_combout ),
	.datad(!\D_ctrl_shift_rot_right~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot_right~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot_right~1 .extended_lut = "off";
defparam \D_ctrl_shift_rot_right~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_ctrl_shift_rot_right~1 .shared_arith = "off";

dffeas R_ctrl_shift_rot_right(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot_right~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_rot_right~q ),
	.prn(vcc));
defparam R_ctrl_shift_rot_right.is_wysiwyg = "true";
defparam R_ctrl_shift_rot_right.power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[3]~13 (
	.dataa(!\E_shift_rot_result[4]~q ),
	.datab(!\E_shift_rot_result[2]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[3]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[3]~13 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[3]~13 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[3]~13 .shared_arith = "off";

dffeas R_ctrl_br(
	.clk(clk_clk),
	.d(\R_ctrl_br_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br~q ),
	.prn(vcc));
defparam R_ctrl_br.is_wysiwyg = "true";
defparam R_ctrl_br.power_up = "low";

cyclonev_lcell_comb \D_ctrl_implicit_dst_eretaddr~2 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_implicit_dst_eretaddr~2 .extended_lut = "off";
defparam \D_ctrl_implicit_dst_eretaddr~2 .lut_mask = 64'h6996966996696996;
defparam \D_ctrl_implicit_dst_eretaddr~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~9 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~9 .extended_lut = "off";
defparam \Equal0~9 .lut_mask = 64'hFFFFFFEFFFFFFFFF;
defparam \Equal0~9 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_retaddr~3 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_retaddr~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_retaddr~3 .extended_lut = "off";
defparam \D_ctrl_retaddr~3 .lut_mask = 64'hF7FFD5FFFFFFFFFF;
defparam \D_ctrl_retaddr~3 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_retaddr~1 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.datac(!\Equal0~9_combout ),
	.datad(!\D_ctrl_exception~1_combout ),
	.datae(!\D_ctrl_retaddr~3_combout ),
	.dataf(!\D_ctrl_retaddr~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_retaddr~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_retaddr~1 .extended_lut = "off";
defparam \D_ctrl_retaddr~1 .lut_mask = 64'hFFFFFFFFFF7FFFFF;
defparam \D_ctrl_retaddr~1 .shared_arith = "off";

dffeas R_ctrl_retaddr(
	.clk(clk_clk),
	.d(\D_ctrl_retaddr~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_retaddr~q ),
	.prn(vcc));
defparam R_ctrl_retaddr.is_wysiwyg = "true";
defparam R_ctrl_retaddr.power_up = "low";

cyclonev_lcell_comb \R_src1~0 (
	.dataa(!\E_valid_from_R~q ),
	.datab(!\R_ctrl_br~q ),
	.datac(!\R_valid~q ),
	.datad(!\R_ctrl_retaddr~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1~0 .extended_lut = "off";
defparam \R_src1~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \R_src1~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_jmp_direct~0 (
	.dataa(!\D_iw[1]~q ),
	.datab(!\D_iw[2]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[4]~q ),
	.datae(!\D_iw[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_jmp_direct~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_jmp_direct~0 .extended_lut = "off";
defparam \D_ctrl_jmp_direct~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \D_ctrl_jmp_direct~0 .shared_arith = "off";

dffeas R_ctrl_jmp_direct(
	.clk(clk_clk),
	.d(\D_ctrl_jmp_direct~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_jmp_direct~q ),
	.prn(vcc));
defparam R_ctrl_jmp_direct.is_wysiwyg = "true";
defparam R_ctrl_jmp_direct.power_up = "low";

cyclonev_lcell_comb \R_src1~1 (
	.dataa(!\E_valid_from_R~q ),
	.datab(!\R_ctrl_jmp_direct~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1~1 .extended_lut = "off";
defparam \R_src1~1 .lut_mask = 64'h7777777777777777;
defparam \R_src1~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h00000000000000FF;
defparam \Add0~57 .shared_arith = "off";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[3]~15 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\Add0~53_sumout ),
	.datad(!\D_iw[7]~q ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[3]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[3]~15 .extended_lut = "off";
defparam \R_src1[3]~15 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[3]~15 .shared_arith = "off";

dffeas \E_src1[3] (
	.clk(clk_clk),
	.d(\R_src1[3]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[3]~q ),
	.prn(vcc));
defparam \E_src1[3] .is_wysiwyg = "true";
defparam \E_src1[3] .power_up = "low";

dffeas \E_shift_rot_result[3] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[3]~13_combout ),
	.asdata(\E_src1[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[3]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[3] .is_wysiwyg = "true";
defparam \E_shift_rot_result[3] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[2]~14 (
	.dataa(!\E_shift_rot_result[3]~q ),
	.datab(!\R_ctrl_shift_rot_right~q ),
	.datac(!\E_shift_rot_result[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[2]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[2]~14 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[2]~14 .lut_mask = 64'h4747474747474747;
defparam \E_shift_rot_result_nxt[2]~14 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[2]~16 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\D_iw[6]~q ),
	.datad(!\Add0~57_sumout ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[2]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[2]~16 .extended_lut = "off";
defparam \R_src1[2]~16 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[2]~16 .shared_arith = "off";

dffeas \E_src1[2] (
	.clk(clk_clk),
	.d(\R_src1[2]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[2]~q ),
	.prn(vcc));
defparam \E_src1[2] .is_wysiwyg = "true";
defparam \E_src1[2] .power_up = "low";

dffeas \E_shift_rot_result[2] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[2]~14_combout ),
	.asdata(\E_src1[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[2]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[2] .is_wysiwyg = "true";
defparam \E_shift_rot_result[2] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[1]~16 (
	.dataa(!\E_shift_rot_result[2]~q ),
	.datab(!\R_ctrl_shift_rot_right~q ),
	.datac(!\E_shift_rot_result[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[1]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[1]~16 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[1]~16 .lut_mask = 64'h4747474747474747;
defparam \E_shift_rot_result_nxt[1]~16 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[26]~0 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[26]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[26]~0 .extended_lut = "off";
defparam \E_src1[26]~0 .lut_mask = 64'h7777777777777777;
defparam \E_src1[26]~0 .shared_arith = "off";

dffeas \E_src1[1] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src1[26]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[1]~q ),
	.prn(vcc));
defparam \E_src1[1] .is_wysiwyg = "true";
defparam \E_src1[1] .power_up = "low";

dffeas \E_shift_rot_result[1] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[1]~16_combout ),
	.asdata(\E_src1[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[1]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[1] .is_wysiwyg = "true";
defparam \E_shift_rot_result[1] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[0]~17 (
	.dataa(!\R_ctrl_shift_rot_right~q ),
	.datab(!\E_shift_rot_result[1]~q ),
	.datac(!\E_shift_rot_fill_bit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[0]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[0]~17 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[0]~17 .lut_mask = 64'h2727272727272727;
defparam \E_shift_rot_result_nxt[0]~17 .shared_arith = "off";

dffeas \E_src1[0] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src1[26]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[0]~q ),
	.prn(vcc));
defparam \E_src1[0] .is_wysiwyg = "true";
defparam \E_src1[0] .power_up = "low";

dffeas \E_shift_rot_result[0] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[0]~17_combout ),
	.asdata(\E_src1[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[0]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[0] .is_wysiwyg = "true";
defparam \E_shift_rot_result[0] .power_up = "low";

cyclonev_lcell_comb \Equal62~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~0 .extended_lut = "off";
defparam \Equal62~0 .lut_mask = 64'hFFFFFFFFFBFFFFFF;
defparam \Equal62~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~2 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~2 .extended_lut = "off";
defparam \Equal62~2 .lut_mask = 64'hFFFFFFFFF7FFFFFF;
defparam \Equal62~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_shift_logical~0 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[15]~q ),
	.datae(!\D_iw[16]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_logical~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_logical~0 .extended_lut = "off";
defparam \D_ctrl_shift_logical~0 .lut_mask = 64'hFFFFFDFFFFFFFDFF;
defparam \D_ctrl_shift_logical~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_shift_logical~1 (
	.dataa(!\Equal62~0_combout ),
	.datab(!\Equal62~2_combout ),
	.datac(!\D_ctrl_shift_logical~0_combout ),
	.datad(!\Equal0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_logical~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_logical~1 .extended_lut = "off";
defparam \D_ctrl_shift_logical~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_ctrl_shift_logical~1 .shared_arith = "off";

dffeas R_ctrl_shift_logical(
	.clk(clk_clk),
	.d(\D_ctrl_shift_logical~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_logical~q ),
	.prn(vcc));
defparam R_ctrl_shift_logical.is_wysiwyg = "true";
defparam R_ctrl_shift_logical.power_up = "low";

cyclonev_lcell_comb \Equal62~1 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~1 .extended_lut = "off";
defparam \Equal62~1 .lut_mask = 64'hFFFFFFFFFFFFF7FF;
defparam \Equal62~1 .shared_arith = "off";

cyclonev_lcell_comb R_ctrl_rot_right_nxt(
	.dataa(!\Equal62~1_combout ),
	.datab(!\Equal0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_ctrl_rot_right_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam R_ctrl_rot_right_nxt.extended_lut = "off";
defparam R_ctrl_rot_right_nxt.lut_mask = 64'h7777777777777777;
defparam R_ctrl_rot_right_nxt.shared_arith = "off";

dffeas R_ctrl_rot_right(
	.clk(clk_clk),
	.d(\R_ctrl_rot_right_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_rot_right~q ),
	.prn(vcc));
defparam R_ctrl_rot_right.is_wysiwyg = "true";
defparam R_ctrl_rot_right.power_up = "low";

cyclonev_lcell_comb \E_shift_rot_fill_bit~0 (
	.dataa(!\E_shift_rot_result[0]~q ),
	.datab(!\R_ctrl_shift_logical~q ),
	.datac(!\R_ctrl_rot_right~q ),
	.datad(!\E_shift_rot_result[31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_fill_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_fill_bit~0 .extended_lut = "off";
defparam \E_shift_rot_fill_bit~0 .lut_mask = 64'hC5FFC5FFC5FFC5FF;
defparam \E_shift_rot_fill_bit~0 .shared_arith = "off";

cyclonev_lcell_comb \E_shift_rot_result_nxt[31]~19 (
	.dataa(!\R_ctrl_shift_rot_right~q ),
	.datab(!\E_shift_rot_fill_bit~0_combout ),
	.datac(!\E_shift_rot_result[30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[31]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[31]~19 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[31]~19 .lut_mask = 64'h2727272727272727;
defparam \E_shift_rot_result_nxt[31]~19 .shared_arith = "off";

dffeas \E_src1[31] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src1[26]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[31]~q ),
	.prn(vcc));
defparam \E_src1[31] .is_wysiwyg = "true";
defparam \E_src1[31] .power_up = "low";

dffeas \E_shift_rot_result[31] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[31]~19_combout ),
	.asdata(\E_src1[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[31]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[31] .is_wysiwyg = "true";
defparam \E_shift_rot_result[31] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[30]~21 (
	.dataa(!\R_ctrl_shift_rot_right~q ),
	.datab(!\E_shift_rot_result[31]~q ),
	.datac(!\E_shift_rot_result[29]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[30]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[30]~21 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[30]~21 .lut_mask = 64'h2727272727272727;
defparam \E_shift_rot_result_nxt[30]~21 .shared_arith = "off";

dffeas \E_src1[30] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src1[26]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[30]~q ),
	.prn(vcc));
defparam \E_src1[30] .is_wysiwyg = "true";
defparam \E_src1[30] .power_up = "low";

dffeas \E_shift_rot_result[30] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[30]~21_combout ),
	.asdata(\E_src1[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[30]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[30] .is_wysiwyg = "true";
defparam \E_shift_rot_result[30] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[29]~31 (
	.dataa(!\R_ctrl_shift_rot_right~q ),
	.datab(!\E_shift_rot_result[30]~q ),
	.datac(!\E_shift_rot_result[28]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[29]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[29]~31 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[29]~31 .lut_mask = 64'h2727272727272727;
defparam \E_shift_rot_result_nxt[29]~31 .shared_arith = "off";

dffeas \E_src1[29] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src1[26]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[29]~q ),
	.prn(vcc));
defparam \E_src1[29] .is_wysiwyg = "true";
defparam \E_src1[29] .power_up = "low";

dffeas \E_shift_rot_result[29] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[29]~31_combout ),
	.asdata(\E_src1[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[29]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[29] .is_wysiwyg = "true";
defparam \E_shift_rot_result[29] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[28]~30 (
	.dataa(!\R_ctrl_shift_rot_right~q ),
	.datab(!\E_shift_rot_result[29]~q ),
	.datac(!\E_shift_rot_result[27]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[28]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[28]~30 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[28]~30 .lut_mask = 64'h2727272727272727;
defparam \E_shift_rot_result_nxt[28]~30 .shared_arith = "off";

dffeas \E_src1[28] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src1[26]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[28]~q ),
	.prn(vcc));
defparam \E_src1[28] .is_wysiwyg = "true";
defparam \E_src1[28] .power_up = "low";

dffeas \E_shift_rot_result[28] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[28]~30_combout ),
	.asdata(\E_src1[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[28]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[28] .is_wysiwyg = "true";
defparam \E_shift_rot_result[28] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[27]~24 (
	.dataa(!\R_ctrl_shift_rot_right~q ),
	.datab(!\E_shift_rot_result[28]~q ),
	.datac(!\E_shift_rot_result[26]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[27]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[27]~24 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[27]~24 .lut_mask = 64'h2727272727272727;
defparam \E_shift_rot_result_nxt[27]~24 .shared_arith = "off";

dffeas \E_src1[27] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src1[26]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[27]~q ),
	.prn(vcc));
defparam \E_src1[27] .is_wysiwyg = "true";
defparam \E_src1[27] .power_up = "low";

dffeas \E_shift_rot_result[27] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[27]~24_combout ),
	.asdata(\E_src1[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[27]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[27] .is_wysiwyg = "true";
defparam \E_shift_rot_result[27] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[26]~29 (
	.dataa(!\R_ctrl_shift_rot_right~q ),
	.datab(!\E_shift_rot_result[25]~q ),
	.datac(!\E_shift_rot_result[27]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[26]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[26]~29 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[26]~29 .lut_mask = 64'h2727272727272727;
defparam \E_shift_rot_result_nxt[26]~29 .shared_arith = "off";

dffeas \E_src1[26] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src1[26]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[26]~q ),
	.prn(vcc));
defparam \E_src1[26] .is_wysiwyg = "true";
defparam \E_src1[26] .power_up = "low";

dffeas \E_shift_rot_result[26] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[26]~29_combout ),
	.asdata(\E_src1[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[26]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[26] .is_wysiwyg = "true";
defparam \E_shift_rot_result[26] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[25]~23 (
	.dataa(!\R_ctrl_shift_rot_right~q ),
	.datab(!\E_shift_rot_result[26]~q ),
	.datac(!\E_shift_rot_result[24]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[25]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[25]~23 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[25]~23 .lut_mask = 64'h2727272727272727;
defparam \E_shift_rot_result_nxt[25]~23 .shared_arith = "off";

dffeas \E_src1[25] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src1[26]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[25]~q ),
	.prn(vcc));
defparam \E_src1[25] .is_wysiwyg = "true";
defparam \E_src1[25] .power_up = "low";

dffeas \E_shift_rot_result[25] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[25]~23_combout ),
	.asdata(\E_src1[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[25]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[25] .is_wysiwyg = "true";
defparam \E_shift_rot_result[25] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[24]~28 (
	.dataa(!\R_ctrl_shift_rot_right~q ),
	.datab(!\E_shift_rot_result[23]~q ),
	.datac(!\E_shift_rot_result[25]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[24]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[24]~28 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[24]~28 .lut_mask = 64'h2727272727272727;
defparam \E_shift_rot_result_nxt[24]~28 .shared_arith = "off";

dffeas \E_src1[24] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src1[26]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[24]~q ),
	.prn(vcc));
defparam \E_src1[24] .is_wysiwyg = "true";
defparam \E_src1[24] .power_up = "low";

dffeas \E_shift_rot_result[24] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[24]~28_combout ),
	.asdata(\E_src1[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[24]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[24] .is_wysiwyg = "true";
defparam \E_shift_rot_result[24] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[23]~27 (
	.dataa(!\R_ctrl_shift_rot_right~q ),
	.datab(!\E_shift_rot_result[22]~q ),
	.datac(!\E_shift_rot_result[24]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[23]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[23]~27 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[23]~27 .lut_mask = 64'h2727272727272727;
defparam \E_shift_rot_result_nxt[23]~27 .shared_arith = "off";

dffeas \E_src1[23] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src1[26]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[23]~q ),
	.prn(vcc));
defparam \E_src1[23] .is_wysiwyg = "true";
defparam \E_src1[23] .power_up = "low";

dffeas \E_shift_rot_result[23] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[23]~27_combout ),
	.asdata(\E_src1[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[23]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[23] .is_wysiwyg = "true";
defparam \E_shift_rot_result[23] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[22]~26 (
	.dataa(!\R_ctrl_shift_rot_right~q ),
	.datab(!\E_shift_rot_result[21]~q ),
	.datac(!\E_shift_rot_result[23]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[22]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[22]~26 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[22]~26 .lut_mask = 64'h2727272727272727;
defparam \E_shift_rot_result_nxt[22]~26 .shared_arith = "off";

dffeas \E_src1[22] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src1[26]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[22]~q ),
	.prn(vcc));
defparam \E_src1[22] .is_wysiwyg = "true";
defparam \E_src1[22] .power_up = "low";

dffeas \E_shift_rot_result[22] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[22]~26_combout ),
	.asdata(\E_src1[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[22]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[22] .is_wysiwyg = "true";
defparam \E_shift_rot_result[22] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[21]~25 (
	.dataa(!\R_ctrl_shift_rot_right~q ),
	.datab(!\E_shift_rot_result[20]~q ),
	.datac(!\E_shift_rot_result[22]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[21]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[21]~25 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[21]~25 .lut_mask = 64'h2727272727272727;
defparam \E_shift_rot_result_nxt[21]~25 .shared_arith = "off";

dffeas \E_src1[21] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src1[26]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[21]~q ),
	.prn(vcc));
defparam \E_src1[21] .is_wysiwyg = "true";
defparam \E_src1[21] .power_up = "low";

dffeas \E_shift_rot_result[21] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[21]~25_combout ),
	.asdata(\E_src1[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[21]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[21] .is_wysiwyg = "true";
defparam \E_shift_rot_result[21] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[20]~22 (
	.dataa(!\R_ctrl_shift_rot_right~q ),
	.datab(!\E_shift_rot_result[19]~q ),
	.datac(!\E_shift_rot_result[21]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[20]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[20]~22 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[20]~22 .lut_mask = 64'h2727272727272727;
defparam \E_shift_rot_result_nxt[20]~22 .shared_arith = "off";

dffeas \E_src1[20] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src1[26]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[20]~q ),
	.prn(vcc));
defparam \E_src1[20] .is_wysiwyg = "true";
defparam \E_src1[20] .power_up = "low";

dffeas \E_shift_rot_result[20] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[20]~22_combout ),
	.asdata(\E_src1[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[20]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[20] .is_wysiwyg = "true";
defparam \E_shift_rot_result[20] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[19]~20 (
	.dataa(!\R_ctrl_shift_rot_right~q ),
	.datab(!\E_shift_rot_result[18]~q ),
	.datac(!\E_shift_rot_result[20]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[19]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[19]~20 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[19]~20 .lut_mask = 64'h2727272727272727;
defparam \E_shift_rot_result_nxt[19]~20 .shared_arith = "off";

dffeas \E_src1[19] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src1[26]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[19]~q ),
	.prn(vcc));
defparam \E_src1[19] .is_wysiwyg = "true";
defparam \E_src1[19] .power_up = "low";

dffeas \E_shift_rot_result[19] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[19]~20_combout ),
	.asdata(\E_src1[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[19]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[19] .is_wysiwyg = "true";
defparam \E_shift_rot_result[19] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[18]~18 (
	.dataa(!\R_ctrl_shift_rot_right~q ),
	.datab(!\E_shift_rot_result[17]~q ),
	.datac(!\E_shift_rot_result[19]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[18]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[18]~18 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[18]~18 .lut_mask = 64'h2727272727272727;
defparam \E_shift_rot_result_nxt[18]~18 .shared_arith = "off";

dffeas \E_src1[18] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src1[26]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[18]~q ),
	.prn(vcc));
defparam \E_src1[18] .is_wysiwyg = "true";
defparam \E_src1[18] .power_up = "low";

dffeas \E_shift_rot_result[18] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[18]~18_combout ),
	.asdata(\E_src1[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[18]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[18] .is_wysiwyg = "true";
defparam \E_shift_rot_result[18] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[17]~15 (
	.dataa(!\E_shift_rot_result[16]~q ),
	.datab(!\R_ctrl_shift_rot_right~q ),
	.datac(!\E_shift_rot_result[18]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[17]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[17]~15 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[17]~15 .lut_mask = 64'h4747474747474747;
defparam \E_shift_rot_result_nxt[17]~15 .shared_arith = "off";

dffeas \E_src1[17] (
	.clk(clk_clk),
	.d(\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src1[26]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[17]~q ),
	.prn(vcc));
defparam \E_src1[17] .is_wysiwyg = "true";
defparam \E_src1[17] .power_up = "low";

dffeas \E_shift_rot_result[17] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[17]~15_combout ),
	.asdata(\E_src1[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[17]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[17] .is_wysiwyg = "true";
defparam \E_shift_rot_result[17] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[16]~12 (
	.dataa(!\E_shift_rot_result[15]~q ),
	.datab(!\R_ctrl_shift_rot_right~q ),
	.datac(!\E_shift_rot_result[17]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[16]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[16]~12 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[16]~12 .lut_mask = 64'h4747474747474747;
defparam \E_shift_rot_result_nxt[16]~12 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[20]~10 (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!av_readdata_pre_201),
	.datad(!q_a_20),
	.datae(!\hbreak_req~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[20]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[20]~10 .extended_lut = "off";
defparam \F_iw[20]~10 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \F_iw[20]~10 .shared_arith = "off";

dffeas \D_iw[20] (
	.clk(clk_clk),
	.d(\F_iw[20]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[20]~q ),
	.prn(vcc));
defparam \D_iw[20] .is_wysiwyg = "true";
defparam \D_iw[20] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000000000FF00;
defparam \Add0~45 .shared_arith = "off";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!F_pc_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[16]~14 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\D_iw[20]~q ),
	.datad(!\Add0~49_sumout ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[16]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[16]~14 .extended_lut = "off";
defparam \R_src1[16]~14 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[16]~14 .shared_arith = "off";

dffeas \E_src1[16] (
	.clk(clk_clk),
	.d(\R_src1[16]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[16]~q ),
	.prn(vcc));
defparam \E_src1[16] .is_wysiwyg = "true";
defparam \E_src1[16] .power_up = "low";

dffeas \E_shift_rot_result[16] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[16]~12_combout ),
	.asdata(\E_src1[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[16]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[16] .is_wysiwyg = "true";
defparam \E_shift_rot_result[16] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[15]~11 (
	.dataa(!\E_shift_rot_result[14]~q ),
	.datab(!\E_shift_rot_result[16]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[15]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[15]~11 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[15]~11 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[15]~11 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[19]~9 (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!av_readdata_pre_191),
	.datad(!q_a_19),
	.datae(!\hbreak_req~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[19]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[19]~9 .extended_lut = "off";
defparam \F_iw[19]~9 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \F_iw[19]~9 .shared_arith = "off";

dffeas \D_iw[19] (
	.clk(clk_clk),
	.d(\F_iw[19]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[19]~q ),
	.prn(vcc));
defparam \D_iw[19] .is_wysiwyg = "true";
defparam \D_iw[19] .power_up = "low";

cyclonev_lcell_comb \R_src1[15]~13 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\D_iw[19]~q ),
	.datad(!\Add0~45_sumout ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[15]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[15]~13 .extended_lut = "off";
defparam \R_src1[15]~13 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[15]~13 .shared_arith = "off";

dffeas \E_src1[15] (
	.clk(clk_clk),
	.d(\R_src1[15]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[15]~q ),
	.prn(vcc));
defparam \E_src1[15] .is_wysiwyg = "true";
defparam \E_src1[15] .power_up = "low";

dffeas \E_shift_rot_result[15] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[15]~11_combout ),
	.asdata(\E_src1[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[15]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[15] .is_wysiwyg = "true";
defparam \E_shift_rot_result[15] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[14]~10 (
	.dataa(!\E_shift_rot_result[13]~q ),
	.datab(!\E_shift_rot_result[15]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[14]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[14]~10 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[14]~10 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[14]~10 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[18]~8 (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!av_readdata_pre_181),
	.datad(!q_a_18),
	.datae(!\hbreak_req~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[18]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[18]~8 .extended_lut = "off";
defparam \F_iw[18]~8 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \F_iw[18]~8 .shared_arith = "off";

dffeas \D_iw[18] (
	.clk(clk_clk),
	.d(\F_iw[18]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[18]~q ),
	.prn(vcc));
defparam \D_iw[18] .is_wysiwyg = "true";
defparam \D_iw[18] .power_up = "low";

cyclonev_lcell_comb \R_src1[14]~12 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\D_iw[18]~q ),
	.datad(!\Add0~41_sumout ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[14]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[14]~12 .extended_lut = "off";
defparam \R_src1[14]~12 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[14]~12 .shared_arith = "off";

dffeas \E_src1[14] (
	.clk(clk_clk),
	.d(\R_src1[14]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[14]~q ),
	.prn(vcc));
defparam \E_src1[14] .is_wysiwyg = "true";
defparam \E_src1[14] .power_up = "low";

dffeas \E_shift_rot_result[14] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[14]~10_combout ),
	.asdata(\E_src1[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[14]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[14] .is_wysiwyg = "true";
defparam \E_shift_rot_result[14] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[13]~9 (
	.dataa(!\E_shift_rot_result[12]~q ),
	.datab(!\E_shift_rot_result[14]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[13]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[13]~9 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[13]~9 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[13]~9 .shared_arith = "off";

dffeas \D_iw[17] (
	.clk(clk_clk),
	.d(src_data_17),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\hbreak_req~0_combout ),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[17]~q ),
	.prn(vcc));
defparam \D_iw[17] .is_wysiwyg = "true";
defparam \D_iw[17] .power_up = "low";

cyclonev_lcell_comb \R_src1[13]~11 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\D_iw[17]~q ),
	.datad(!\Add0~37_sumout ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[13]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[13]~11 .extended_lut = "off";
defparam \R_src1[13]~11 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[13]~11 .shared_arith = "off";

dffeas \E_src1[13] (
	.clk(clk_clk),
	.d(\R_src1[13]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[13]~q ),
	.prn(vcc));
defparam \E_src1[13] .is_wysiwyg = "true";
defparam \E_src1[13] .power_up = "low";

dffeas \E_shift_rot_result[13] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[13]~9_combout ),
	.asdata(\E_src1[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[13]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[13] .is_wysiwyg = "true";
defparam \E_shift_rot_result[13] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[12]~8 (
	.dataa(!\E_shift_rot_result[11]~q ),
	.datab(!\E_shift_rot_result[13]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[12]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[12]~8 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[12]~8 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[12]~8 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[12]~10 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\R_src1~0_combout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\Add0~33_sumout ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[12]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[12]~10 .extended_lut = "off";
defparam \R_src1[12]~10 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src1[12]~10 .shared_arith = "off";

dffeas \E_src1[12] (
	.clk(clk_clk),
	.d(\R_src1[12]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[12]~q ),
	.prn(vcc));
defparam \E_src1[12] .is_wysiwyg = "true";
defparam \E_src1[12] .power_up = "low";

dffeas \E_shift_rot_result[12] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[12]~8_combout ),
	.asdata(\E_src1[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[12]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[12] .is_wysiwyg = "true";
defparam \E_shift_rot_result[12] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[11]~1 (
	.dataa(!\E_shift_rot_result[10]~q ),
	.datab(!\E_shift_rot_result[12]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[11]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[11]~1 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[11]~1 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[11]~1 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[11]~3 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\R_src1~0_combout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\Add0~5_sumout ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[11]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[11]~3 .extended_lut = "off";
defparam \R_src1[11]~3 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src1[11]~3 .shared_arith = "off";

dffeas \E_src1[11] (
	.clk(clk_clk),
	.d(\R_src1[11]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[11]~q ),
	.prn(vcc));
defparam \E_src1[11] .is_wysiwyg = "true";
defparam \E_src1[11] .power_up = "low";

dffeas \E_shift_rot_result[11] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[11]~1_combout ),
	.asdata(\E_src1[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[11]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[11] .is_wysiwyg = "true";
defparam \E_shift_rot_result[11] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[10]~2 (
	.dataa(!\E_shift_rot_result[11]~q ),
	.datab(!\E_shift_rot_result[9]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[10]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[10]~2 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[10]~2 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[10]~2 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[10]~4 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\R_src1~0_combout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\Add0~9_sumout ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[10]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[10]~4 .extended_lut = "off";
defparam \R_src1[10]~4 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src1[10]~4 .shared_arith = "off";

dffeas \E_src1[10] (
	.clk(clk_clk),
	.d(\R_src1[10]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[10]~q ),
	.prn(vcc));
defparam \E_src1[10] .is_wysiwyg = "true";
defparam \E_src1[10] .power_up = "low";

dffeas \E_shift_rot_result[10] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[10]~2_combout ),
	.asdata(\E_src1[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[10]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[10] .is_wysiwyg = "true";
defparam \E_shift_rot_result[10] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[9]~3 (
	.dataa(!\E_shift_rot_result[10]~q ),
	.datab(!\E_shift_rot_result[8]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[9]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[9]~3 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[9]~3 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[9]~3 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[9]~5 (
	.dataa(!\D_iw[13]~q ),
	.datab(!\R_src1~0_combout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\Add0~13_sumout ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[9]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[9]~5 .extended_lut = "off";
defparam \R_src1[9]~5 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src1[9]~5 .shared_arith = "off";

dffeas \E_src1[9] (
	.clk(clk_clk),
	.d(\R_src1[9]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[9]~q ),
	.prn(vcc));
defparam \E_src1[9] .is_wysiwyg = "true";
defparam \E_src1[9] .power_up = "low";

dffeas \E_shift_rot_result[9] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[9]~3_combout ),
	.asdata(\E_src1[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[9]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[9] .is_wysiwyg = "true";
defparam \E_shift_rot_result[9] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[8]~4 (
	.dataa(!\E_shift_rot_result[9]~q ),
	.datab(!\E_shift_rot_result[7]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[8]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[8]~4 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[8]~4 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[8]~4 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[8]~6 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\R_src1~0_combout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\Add0~17_sumout ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[8]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[8]~6 .extended_lut = "off";
defparam \R_src1[8]~6 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src1[8]~6 .shared_arith = "off";

dffeas \E_src1[8] (
	.clk(clk_clk),
	.d(\R_src1[8]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[8]~q ),
	.prn(vcc));
defparam \E_src1[8] .is_wysiwyg = "true";
defparam \E_src1[8] .power_up = "low";

dffeas \E_shift_rot_result[8] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[8]~4_combout ),
	.asdata(\E_src1[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[8]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[8] .is_wysiwyg = "true";
defparam \E_shift_rot_result[8] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[7]~5 (
	.dataa(!\E_shift_rot_result[8]~q ),
	.datab(!\E_shift_rot_result[6]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[7]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[7]~5 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[7]~5 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[7]~5 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[7]~7 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\R_src1~0_combout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\Add0~21_sumout ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[7]~7 .extended_lut = "off";
defparam \R_src1[7]~7 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src1[7]~7 .shared_arith = "off";

dffeas \E_src1[7] (
	.clk(clk_clk),
	.d(\R_src1[7]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[7]~q ),
	.prn(vcc));
defparam \E_src1[7] .is_wysiwyg = "true";
defparam \E_src1[7] .power_up = "low";

dffeas \E_shift_rot_result[7] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[7]~5_combout ),
	.asdata(\E_src1[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[7]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[7] .is_wysiwyg = "true";
defparam \E_shift_rot_result[7] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[6]~6 (
	.dataa(!\E_shift_rot_result[7]~q ),
	.datab(!\E_shift_rot_result[5]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[6]~6 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[6]~6 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[6]~8 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\D_iw[10]~q ),
	.datad(!\Add0~25_sumout ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[6]~8 .extended_lut = "off";
defparam \R_src1[6]~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[6]~8 .shared_arith = "off";

dffeas \E_src1[6] (
	.clk(clk_clk),
	.d(\R_src1[6]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[6]~q ),
	.prn(vcc));
defparam \E_src1[6] .is_wysiwyg = "true";
defparam \E_src1[6] .power_up = "low";

dffeas \E_shift_rot_result[6] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[6]~6_combout ),
	.asdata(\E_src1[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[6]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[6] .is_wysiwyg = "true";
defparam \E_shift_rot_result[6] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[5]~7 (
	.dataa(!\E_shift_rot_result[4]~q ),
	.datab(!\E_shift_rot_result[6]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[5]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[5]~7 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[5]~7 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[5]~7 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[5]~9 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\R_src1~1_combout ),
	.datac(!\Add0~29_sumout ),
	.datad(!\D_iw[9]~q ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[5]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[5]~9 .extended_lut = "off";
defparam \R_src1[5]~9 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src1[5]~9 .shared_arith = "off";

dffeas \E_src1[5] (
	.clk(clk_clk),
	.d(\R_src1[5]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[5]~q ),
	.prn(vcc));
defparam \E_src1[5] .is_wysiwyg = "true";
defparam \E_src1[5] .power_up = "low";

dffeas \E_shift_rot_result[5] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[5]~7_combout ),
	.asdata(\E_src1[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[5]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[5] .is_wysiwyg = "true";
defparam \E_shift_rot_result[5] .power_up = "low";

cyclonev_lcell_comb \E_shift_rot_result_nxt[4]~0 (
	.dataa(!\E_shift_rot_result[5]~q ),
	.datab(!\E_shift_rot_result[3]~q ),
	.datac(!\R_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_shift_rot_result_nxt[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_shift_rot_result_nxt[4]~0 .extended_lut = "off";
defparam \E_shift_rot_result_nxt[4]~0 .lut_mask = 64'h5353535353535353;
defparam \E_shift_rot_result_nxt[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \R_src1[4]~2 (
	.dataa(!\R_src1~0_combout ),
	.datab(!\Add0~1_sumout ),
	.datac(!\R_src1~1_combout ),
	.datad(!\D_iw[8]~q ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src1[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src1[4]~2 .extended_lut = "off";
defparam \R_src1[4]~2 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \R_src1[4]~2 .shared_arith = "off";

dffeas \E_src1[4] (
	.clk(clk_clk),
	.d(\R_src1[4]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[4]~q ),
	.prn(vcc));
defparam \E_src1[4] .is_wysiwyg = "true";
defparam \E_src1[4] .power_up = "low";

dffeas \E_shift_rot_result[4] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[4]~0_combout ),
	.asdata(\E_src1[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[4]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[4] .is_wysiwyg = "true";
defparam \E_shift_rot_result[4] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_logic~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[16]~q ),
	.datae(!\Equal0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_logic~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_logic~0 .extended_lut = "off";
defparam \D_ctrl_logic~0 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \D_ctrl_logic~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_logic~1 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[0]~q ),
	.dataf(!\D_ctrl_logic~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_logic~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_logic~1 .extended_lut = "off";
defparam \D_ctrl_logic~1 .lut_mask = 64'hFFFFFF7FFFFFFFFF;
defparam \D_ctrl_logic~1 .shared_arith = "off";

dffeas R_ctrl_logic(
	.clk(clk_clk),
	.d(\D_ctrl_logic~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_logic~q ),
	.prn(vcc));
defparam R_ctrl_logic.is_wysiwyg = "true";
defparam R_ctrl_logic.power_up = "low";

cyclonev_lcell_comb \D_logic_op_raw[1]~0 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\Equal0~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op_raw[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op_raw[1]~0 .extended_lut = "off";
defparam \D_logic_op_raw[1]~0 .lut_mask = 64'h5353535353535353;
defparam \D_logic_op_raw[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_force_xor~1 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_force_xor~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_force_xor~1 .extended_lut = "off";
defparam \D_ctrl_alu_force_xor~1 .lut_mask = 64'hFFFFFFFFFFFFDF8F;
defparam \D_ctrl_alu_force_xor~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_subtract~2 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_subtract~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_subtract~2 .extended_lut = "off";
defparam \D_ctrl_alu_subtract~2 .lut_mask = 64'hFFFFBFFBFFFFBFFB;
defparam \D_ctrl_alu_subtract~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_force_xor~0 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_force_xor~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_force_xor~0 .extended_lut = "off";
defparam \D_ctrl_alu_force_xor~0 .lut_mask = 64'hFFFFFFFF96696996;
defparam \D_ctrl_alu_force_xor~0 .shared_arith = "off";

cyclonev_lcell_comb \D_logic_op[1]~0 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\D_logic_op_raw[1]~0_combout ),
	.datac(!\D_ctrl_alu_force_xor~1_combout ),
	.datad(!\D_ctrl_alu_subtract~2_combout ),
	.datae(!\D_ctrl_alu_force_xor~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op[1]~0 .extended_lut = "off";
defparam \D_logic_op[1]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \D_logic_op[1]~0 .shared_arith = "off";

dffeas \R_logic_op[1] (
	.clk(clk_clk),
	.d(\D_logic_op[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_logic_op[1]~q ),
	.prn(vcc));
defparam \R_logic_op[1] .is_wysiwyg = "true";
defparam \R_logic_op[1] .power_up = "low";

cyclonev_lcell_comb \D_logic_op_raw[0]~1 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\Equal0~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op_raw[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op_raw[0]~1 .extended_lut = "off";
defparam \D_logic_op_raw[0]~1 .lut_mask = 64'h5353535353535353;
defparam \D_logic_op_raw[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \D_logic_op[0]~1 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\D_ctrl_alu_force_xor~1_combout ),
	.datac(!\D_ctrl_alu_subtract~2_combout ),
	.datad(!\D_ctrl_alu_force_xor~0_combout ),
	.datae(!\D_logic_op_raw[0]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op[0]~1 .extended_lut = "off";
defparam \D_logic_op[0]~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \D_logic_op[0]~1 .shared_arith = "off";

dffeas \R_logic_op[0] (
	.clk(clk_clk),
	.d(\D_logic_op[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_logic_op[0]~q ),
	.prn(vcc));
defparam \R_logic_op[0] .is_wysiwyg = "true";
defparam \R_logic_op[0] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[4]~0 (
	.dataa(!\E_src1[4]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\R_logic_op[1]~q ),
	.datad(!\R_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[4]~0 .extended_lut = "off";
defparam \E_logic_result[4]~0 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_subtract~1 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_subtract~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_subtract~1 .extended_lut = "off";
defparam \D_ctrl_alu_subtract~1 .lut_mask = 64'hFFFFFFD7FFFFFF7D;
defparam \D_ctrl_alu_subtract~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_subtract~0 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_subtract~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_subtract~0 .extended_lut = "off";
defparam \D_ctrl_alu_subtract~0 .lut_mask = 64'hFFFFDFFDFFFFDFFD;
defparam \D_ctrl_alu_subtract~0 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_sub~0 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\R_valid~q ),
	.datac(!\D_ctrl_alu_subtract~2_combout ),
	.datad(!\D_ctrl_alu_subtract~1_combout ),
	.datae(!\D_ctrl_alu_subtract~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_sub~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_sub~0 .extended_lut = "off";
defparam \E_alu_sub~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_sub~0 .shared_arith = "off";

dffeas E_alu_sub(
	.clk(clk_clk),
	.d(\E_alu_sub~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_alu_sub~q ),
	.prn(vcc));
defparam E_alu_sub.is_wysiwyg = "true";
defparam E_alu_sub.power_up = "low";

cyclonev_lcell_comb \Add2~78 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add2~78_cout ),
	.shareout());
defparam \Add2~78 .extended_lut = "off";
defparam \Add2~78 .lut_mask = 64'h0000000000005555;
defparam \Add2~78 .shared_arith = "off";

cyclonev_lcell_comb \Add2~69 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[0]~q ),
	.datae(gnd),
	.dataf(!\E_src1[0]~q ),
	.datag(gnd),
	.cin(\Add2~78_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~69_sumout ),
	.cout(\Add2~70 ),
	.shareout());
defparam \Add2~69 .extended_lut = "off";
defparam \Add2~69 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~69 .shared_arith = "off";

cyclonev_lcell_comb \Add2~61 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[1]~q ),
	.datae(gnd),
	.dataf(!\E_src1[1]~q ),
	.datag(gnd),
	.cin(\Add2~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~61_sumout ),
	.cout(\Add2~62 ),
	.shareout());
defparam \Add2~61 .extended_lut = "off";
defparam \Add2~61 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~61 .shared_arith = "off";

cyclonev_lcell_comb \Add2~57 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[2]~q ),
	.datae(gnd),
	.dataf(!\E_src1[2]~q ),
	.datag(gnd),
	.cin(\Add2~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~57_sumout ),
	.cout(\Add2~58 ),
	.shareout());
defparam \Add2~57 .extended_lut = "off";
defparam \Add2~57 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~57 .shared_arith = "off";

cyclonev_lcell_comb \Add2~53 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[3]~q ),
	.datae(gnd),
	.dataf(!\E_src1[3]~q ),
	.datag(gnd),
	.cin(\Add2~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~53_sumout ),
	.cout(\Add2~54 ),
	.shareout());
defparam \Add2~53 .extended_lut = "off";
defparam \Add2~53 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~53 .shared_arith = "off";

cyclonev_lcell_comb \Add2~1 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[4]~q ),
	.datae(gnd),
	.dataf(!\E_src1[4]~q ),
	.datag(gnd),
	.cin(\Add2~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~1_sumout ),
	.cout(\Add2~2 ),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~1 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[4]~0 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\E_shift_rot_result[4]~q ),
	.datac(!\R_ctrl_logic~q ),
	.datad(!\E_logic_result[4]~0_combout ),
	.datae(!\Add2~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[4]~0 .extended_lut = "off";
defparam \E_alu_result[4]~0 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \E_alu_result[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~4 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~4 .extended_lut = "off";
defparam \Equal62~4 .lut_mask = 64'hFFFFFFBFFFFFFFFF;
defparam \Equal62~4 .shared_arith = "off";

cyclonev_lcell_comb D_op_rdctl(
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal62~4_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_op_rdctl~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_op_rdctl.extended_lut = "off";
defparam D_op_rdctl.lut_mask = 64'h7777777777777777;
defparam D_op_rdctl.shared_arith = "off";

dffeas R_ctrl_rd_ctl_reg(
	.clk(clk_clk),
	.d(\D_op_rdctl~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_rd_ctl_reg~q ),
	.prn(vcc));
defparam R_ctrl_rd_ctl_reg.is_wysiwyg = "true";
defparam R_ctrl_rd_ctl_reg.power_up = "low";

cyclonev_lcell_comb \Equal62~5 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~5 .extended_lut = "off";
defparam \Equal62~5 .lut_mask = 64'hFFFFFFFFFFFEFFFF;
defparam \Equal62~5 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~6 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~6 .extended_lut = "off";
defparam \Equal62~6 .lut_mask = 64'hFFFEFFFFFFFFFFFF;
defparam \Equal62~6 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_unsigned_lo_imm16~1 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_unsigned_lo_imm16~1 .extended_lut = "off";
defparam \D_ctrl_unsigned_lo_imm16~1 .lut_mask = 64'hFFFFFFFFFFFFFF7D;
defparam \D_ctrl_unsigned_lo_imm16~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'hFFFFFFFFFFFFFEFF;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~4 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~4 .extended_lut = "off";
defparam \Equal0~4 .lut_mask = 64'hFFFFFFFFFEFFFFFF;
defparam \Equal0~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~5 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~5 .extended_lut = "off";
defparam \Equal0~5 .lut_mask = 64'hFFFFFFFEFFFFFFFF;
defparam \Equal0~5 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~6 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~6 .extended_lut = "off";
defparam \Equal0~6 .lut_mask = 64'hFFFFFFFFFFFEFFFF;
defparam \Equal0~6 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_br_cmp~0 (
	.dataa(!\Equal0~1_combout ),
	.datab(!\Equal0~4_combout ),
	.datac(!\Equal0~5_combout ),
	.datad(!\Equal0~6_combout ),
	.datae(!\R_ctrl_br_nxt~0_combout ),
	.dataf(!\R_ctrl_br_nxt~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_br_cmp~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_br_cmp~0 .extended_lut = "off";
defparam \D_ctrl_br_cmp~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \D_ctrl_br_cmp~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_br_cmp~1 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\D_ctrl_alu_force_xor~1_combout ),
	.datac(!\Equal62~5_combout ),
	.datad(!\Equal62~6_combout ),
	.datae(!\D_ctrl_unsigned_lo_imm16~1_combout ),
	.dataf(!\D_ctrl_br_cmp~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_br_cmp~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_br_cmp~1 .extended_lut = "off";
defparam \D_ctrl_br_cmp~1 .lut_mask = 64'hFFFFFFFF7FFFFFFF;
defparam \D_ctrl_br_cmp~1 .shared_arith = "off";

dffeas R_ctrl_br_cmp(
	.clk(clk_clk),
	.d(\D_ctrl_br_cmp~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br_cmp~q ),
	.prn(vcc));
defparam R_ctrl_br_cmp.is_wysiwyg = "true";
defparam R_ctrl_br_cmp.power_up = "low";

cyclonev_lcell_comb \E_alu_result~1 (
	.dataa(!\R_ctrl_rd_ctl_reg~q ),
	.datab(!\R_ctrl_br_cmp~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~1 .extended_lut = "off";
defparam \E_alu_result~1 .lut_mask = 64'h7777777777777777;
defparam \E_alu_result~1 .shared_arith = "off";

cyclonev_lcell_comb \E_src2[15]~0 (
	.dataa(!\R_ctrl_src_imm5_shift_rot~q ),
	.datab(!\R_ctrl_hi_imm16~q ),
	.datac(!\R_ctrl_force_src2_zero~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src2[15]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src2[15]~0 .extended_lut = "off";
defparam \E_src2[15]~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_src2[15]~0 .shared_arith = "off";

dffeas \E_src2[11] (
	.clk(clk_clk),
	.d(\D_iw[17]~q ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[15]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[11]~q ),
	.prn(vcc));
defparam \E_src2[11] .is_wysiwyg = "true";
defparam \E_src2[11] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[11]~1 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[11]~q ),
	.datad(!\E_src2[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[11]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[11]~1 .extended_lut = "off";
defparam \E_logic_result[11]~1 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[11]~1 .shared_arith = "off";

dffeas \E_src2[10] (
	.clk(clk_clk),
	.d(\D_iw[16]~q ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[15]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[10]~q ),
	.prn(vcc));
defparam \E_src2[10] .is_wysiwyg = "true";
defparam \E_src2[10] .power_up = "low";

dffeas \E_src2[9] (
	.clk(clk_clk),
	.d(\D_iw[15]~q ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[15]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[9]~q ),
	.prn(vcc));
defparam \E_src2[9] .is_wysiwyg = "true";
defparam \E_src2[9] .power_up = "low";

dffeas \E_src2[8] (
	.clk(clk_clk),
	.d(\D_iw[14]~q ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[15]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[8]~q ),
	.prn(vcc));
defparam \E_src2[8] .is_wysiwyg = "true";
defparam \E_src2[8] .power_up = "low";

dffeas \E_src2[7] (
	.clk(clk_clk),
	.d(\D_iw[13]~q ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[15]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[7]~q ),
	.prn(vcc));
defparam \E_src2[7] .is_wysiwyg = "true";
defparam \E_src2[7] .power_up = "low";

dffeas \E_src2[6] (
	.clk(clk_clk),
	.d(\D_iw[12]~q ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[15]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[6]~q ),
	.prn(vcc));
defparam \E_src2[6] .is_wysiwyg = "true";
defparam \E_src2[6] .power_up = "low";

dffeas \E_src2[5] (
	.clk(clk_clk),
	.d(\D_iw[11]~q ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[15]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[5]~q ),
	.prn(vcc));
defparam \E_src2[5] .is_wysiwyg = "true";
defparam \E_src2[5] .power_up = "low";

cyclonev_lcell_comb \Add2~29 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[5]~q ),
	.datae(gnd),
	.dataf(!\E_src1[5]~q ),
	.datag(gnd),
	.cin(\Add2~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~29_sumout ),
	.cout(\Add2~30 ),
	.shareout());
defparam \Add2~29 .extended_lut = "off";
defparam \Add2~29 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~29 .shared_arith = "off";

cyclonev_lcell_comb \Add2~25 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[6]~q ),
	.datae(gnd),
	.dataf(!\E_src1[6]~q ),
	.datag(gnd),
	.cin(\Add2~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~25_sumout ),
	.cout(\Add2~26 ),
	.shareout());
defparam \Add2~25 .extended_lut = "off";
defparam \Add2~25 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~25 .shared_arith = "off";

cyclonev_lcell_comb \Add2~21 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[7]~q ),
	.datae(gnd),
	.dataf(!\E_src1[7]~q ),
	.datag(gnd),
	.cin(\Add2~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~21_sumout ),
	.cout(\Add2~22 ),
	.shareout());
defparam \Add2~21 .extended_lut = "off";
defparam \Add2~21 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~21 .shared_arith = "off";

cyclonev_lcell_comb \Add2~17 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[8]~q ),
	.datae(gnd),
	.dataf(!\E_src1[8]~q ),
	.datag(gnd),
	.cin(\Add2~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~17_sumout ),
	.cout(\Add2~18 ),
	.shareout());
defparam \Add2~17 .extended_lut = "off";
defparam \Add2~17 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~17 .shared_arith = "off";

cyclonev_lcell_comb \Add2~13 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[9]~q ),
	.datae(gnd),
	.dataf(!\E_src1[9]~q ),
	.datag(gnd),
	.cin(\Add2~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~13_sumout ),
	.cout(\Add2~14 ),
	.shareout());
defparam \Add2~13 .extended_lut = "off";
defparam \Add2~13 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~13 .shared_arith = "off";

cyclonev_lcell_comb \Add2~9 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[10]~q ),
	.datae(gnd),
	.dataf(!\E_src1[10]~q ),
	.datag(gnd),
	.cin(\Add2~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~9_sumout ),
	.cout(\Add2~10 ),
	.shareout());
defparam \Add2~9 .extended_lut = "off";
defparam \Add2~9 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~9 .shared_arith = "off";

cyclonev_lcell_comb \Add2~5 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[11]~q ),
	.datae(gnd),
	.dataf(!\E_src1[11]~q ),
	.datag(gnd),
	.cin(\Add2~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~5_sumout ),
	.cout(\Add2~6 ),
	.shareout());
defparam \Add2~5 .extended_lut = "off";
defparam \Add2~5 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~5 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[11]~2 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[11]~q ),
	.datad(!\E_logic_result[11]~1_combout ),
	.datae(!\Add2~5_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[11]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[11]~2 .extended_lut = "off";
defparam \E_alu_result[11]~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[11]~2 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[10]~2 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[10]~q ),
	.datad(!\E_src1[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[10]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[10]~2 .extended_lut = "off";
defparam \E_logic_result[10]~2 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[10]~2 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[10]~3 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[10]~q ),
	.datad(!\E_logic_result[10]~2_combout ),
	.datae(!\Add2~9_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[10]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[10]~3 .extended_lut = "off";
defparam \E_alu_result[10]~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[10]~3 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[9]~3 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[9]~q ),
	.datad(!\E_src1[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[9]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[9]~3 .extended_lut = "off";
defparam \E_logic_result[9]~3 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[9]~3 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[9]~4 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[9]~q ),
	.datad(!\E_logic_result[9]~3_combout ),
	.datae(!\Add2~13_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[9]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[9]~4 .extended_lut = "off";
defparam \E_alu_result[9]~4 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[9]~4 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[8]~4 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[8]~q ),
	.datad(!\E_src1[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[8]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[8]~4 .extended_lut = "off";
defparam \E_logic_result[8]~4 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[8]~4 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[8]~5 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[8]~q ),
	.datad(!\E_logic_result[8]~4_combout ),
	.datae(!\Add2~17_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[8]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[8]~5 .extended_lut = "off";
defparam \E_alu_result[8]~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[8]~5 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[7]~5 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[7]~q ),
	.datad(!\E_src1[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[7]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[7]~5 .extended_lut = "off";
defparam \E_logic_result[7]~5 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[7]~5 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[7]~6 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[7]~q ),
	.datad(!\E_logic_result[7]~5_combout ),
	.datae(!\Add2~21_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[7]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[7]~6 .extended_lut = "off";
defparam \E_alu_result[7]~6 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[7]~6 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[6]~6 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[6]~q ),
	.datad(!\E_src1[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[6]~6 .extended_lut = "off";
defparam \E_logic_result[6]~6 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[6]~7 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[6]~q ),
	.datad(!\E_logic_result[6]~6_combout ),
	.datae(!\Add2~25_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[6]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[6]~7 .extended_lut = "off";
defparam \E_alu_result[6]~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[6]~7 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[5]~7 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[5]~q ),
	.datad(!\E_src1[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[5]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[5]~7 .extended_lut = "off";
defparam \E_logic_result[5]~7 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[5]~7 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[5]~8 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[5]~q ),
	.datad(!\E_logic_result[5]~7_combout ),
	.datae(!\Add2~29_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[5]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[5]~8 .extended_lut = "off";
defparam \E_alu_result[5]~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[5]~8 .shared_arith = "off";

dffeas \E_src2[12] (
	.clk(clk_clk),
	.d(\D_iw[18]~q ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[15]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[12]~q ),
	.prn(vcc));
defparam \E_src2[12] .is_wysiwyg = "true";
defparam \E_src2[12] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[12]~8 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[12]~q ),
	.datad(!\E_src2[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[12]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[12]~8 .extended_lut = "off";
defparam \E_logic_result[12]~8 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[12]~8 .shared_arith = "off";

cyclonev_lcell_comb \Add2~33 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[12]~q ),
	.datae(gnd),
	.dataf(!\E_src1[12]~q ),
	.datag(gnd),
	.cin(\Add2~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~33_sumout ),
	.cout(\Add2~34 ),
	.shareout());
defparam \Add2~33 .extended_lut = "off";
defparam \Add2~33 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~33 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[12]~9 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[12]~q ),
	.datad(!\E_logic_result[12]~8_combout ),
	.datae(!\Add2~33_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[12]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[12]~9 .extended_lut = "off";
defparam \E_alu_result[12]~9 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[12]~9 .shared_arith = "off";

dffeas \E_src2[13] (
	.clk(clk_clk),
	.d(\D_iw[19]~q ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[15]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[13]~q ),
	.prn(vcc));
defparam \E_src2[13] .is_wysiwyg = "true";
defparam \E_src2[13] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[13]~9 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[13]~q ),
	.datad(!\E_src2[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[13]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[13]~9 .extended_lut = "off";
defparam \E_logic_result[13]~9 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[13]~9 .shared_arith = "off";

cyclonev_lcell_comb \Add2~37 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[13]~q ),
	.datae(gnd),
	.dataf(!\E_src1[13]~q ),
	.datag(gnd),
	.cin(\Add2~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~37_sumout ),
	.cout(\Add2~38 ),
	.shareout());
defparam \Add2~37 .extended_lut = "off";
defparam \Add2~37 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~37 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[13]~10 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[13]~q ),
	.datad(!\E_logic_result[13]~9_combout ),
	.datae(!\Add2~37_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[13]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[13]~10 .extended_lut = "off";
defparam \E_alu_result[13]~10 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[13]~10 .shared_arith = "off";

dffeas \E_src2[14] (
	.clk(clk_clk),
	.d(\D_iw[20]~q ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[15]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[14]~q ),
	.prn(vcc));
defparam \E_src2[14] .is_wysiwyg = "true";
defparam \E_src2[14] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[14]~10 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[14]~q ),
	.datad(!\E_src2[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[14]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[14]~10 .extended_lut = "off";
defparam \E_logic_result[14]~10 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[14]~10 .shared_arith = "off";

cyclonev_lcell_comb \Add2~41 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[14]~q ),
	.datae(gnd),
	.dataf(!\E_src1[14]~q ),
	.datag(gnd),
	.cin(\Add2~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~41_sumout ),
	.cout(\Add2~42 ),
	.shareout());
defparam \Add2~41 .extended_lut = "off";
defparam \Add2~41 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~41 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[14]~11 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[14]~q ),
	.datad(!\E_logic_result[14]~10_combout ),
	.datae(!\Add2~41_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[14]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[14]~11 .extended_lut = "off";
defparam \E_alu_result[14]~11 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[14]~11 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[21]~11 (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!av_readdata_pre_211),
	.datad(!q_a_21),
	.datae(!\hbreak_req~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[21]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[21]~11 .extended_lut = "off";
defparam \F_iw[21]~11 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \F_iw[21]~11 .shared_arith = "off";

dffeas \D_iw[21] (
	.clk(clk_clk),
	.d(\F_iw[21]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[21]~q ),
	.prn(vcc));
defparam \D_iw[21] .is_wysiwyg = "true";
defparam \D_iw[21] .power_up = "low";

dffeas \E_src2[15] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_src2[15]~0_combout ),
	.sload(!\R_src2_use_imm~q ),
	.ena(vcc),
	.q(\E_src2[15]~q ),
	.prn(vcc));
defparam \E_src2[15] .is_wysiwyg = "true";
defparam \E_src2[15] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[15]~11 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[15]~q ),
	.datad(!\E_src2[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[15]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[15]~11 .extended_lut = "off";
defparam \E_logic_result[15]~11 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[15]~11 .shared_arith = "off";

cyclonev_lcell_comb \Add2~45 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[15]~q ),
	.datae(gnd),
	.dataf(!\E_src1[15]~q ),
	.datag(gnd),
	.cin(\Add2~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~45_sumout ),
	.cout(\Add2~46 ),
	.shareout());
defparam \Add2~45 .extended_lut = "off";
defparam \Add2~45 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~45 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[15]~12 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[15]~q ),
	.datad(!\E_logic_result[15]~11_combout ),
	.datae(!\Add2~45_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[15]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[15]~12 .extended_lut = "off";
defparam \E_alu_result[15]~12 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[15]~12 .shared_arith = "off";

cyclonev_lcell_comb \R_src2_hi[0]~0 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\R_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_iw[6]~q ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[0]~0 .extended_lut = "off";
defparam \R_src2_hi[0]~0 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src2_hi[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_logic~2 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_logic~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_logic~2 .extended_lut = "off";
defparam \D_ctrl_logic~2 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \D_ctrl_logic~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_unsigned_lo_imm16~0 (
	.dataa(!\D_ctrl_unsigned_lo_imm16~1_combout ),
	.datab(!\R_src2_use_imm~1_combout ),
	.datac(!\D_ctrl_logic~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_unsigned_lo_imm16~0 .extended_lut = "off";
defparam \D_ctrl_unsigned_lo_imm16~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \D_ctrl_unsigned_lo_imm16~0 .shared_arith = "off";

dffeas R_ctrl_unsigned_lo_imm16(
	.clk(clk_clk),
	.d(\D_ctrl_unsigned_lo_imm16~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_unsigned_lo_imm16~q ),
	.prn(vcc));
defparam R_ctrl_unsigned_lo_imm16.is_wysiwyg = "true";
defparam R_ctrl_unsigned_lo_imm16.power_up = "low";

cyclonev_lcell_comb \R_src2_hi~1 (
	.dataa(!\R_ctrl_force_src2_zero~q ),
	.datab(!\R_ctrl_unsigned_lo_imm16~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi~1 .extended_lut = "off";
defparam \R_src2_hi~1 .lut_mask = 64'h7777777777777777;
defparam \R_src2_hi~1 .shared_arith = "off";

dffeas \E_src2[16] (
	.clk(clk_clk),
	.d(\R_src2_hi[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[16]~q ),
	.prn(vcc));
defparam \E_src2[16] .is_wysiwyg = "true";
defparam \E_src2[16] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[16]~12 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[16]~q ),
	.datad(!\E_src2[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[16]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[16]~12 .extended_lut = "off";
defparam \E_logic_result[16]~12 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[16]~12 .shared_arith = "off";

cyclonev_lcell_comb \Add2~49 (
	.dataa(!\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[16]~q ),
	.datae(gnd),
	.dataf(!\E_src1[16]~q ),
	.datag(gnd),
	.cin(\Add2~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~49_sumout ),
	.cout(\Add2~50 ),
	.shareout());
defparam \Add2~49 .extended_lut = "off";
defparam \Add2~49 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~49 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[16]~13 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[16]~q ),
	.datad(!\E_logic_result[16]~12_combout ),
	.datae(!\Add2~49_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[16]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[16]~13 .extended_lut = "off";
defparam \E_alu_result[16]~13 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[16]~13 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[3]~13 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[3]~q ),
	.datad(!\E_src1[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[3]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[3]~13 .extended_lut = "off";
defparam \E_logic_result[3]~13 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[3]~13 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[3]~14 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[3]~q ),
	.datad(!\E_logic_result[3]~13_combout ),
	.datae(!\Add2~53_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[3]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[3]~14 .extended_lut = "off";
defparam \E_alu_result[3]~14 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[3]~14 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[2]~14 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[2]~q ),
	.datad(!\E_src1[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[2]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[2]~14 .extended_lut = "off";
defparam \E_logic_result[2]~14 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[2]~14 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[2]~15 (
	.dataa(!\R_ctrl_shift_rot~q ),
	.datab(!\R_ctrl_logic~q ),
	.datac(!\E_shift_rot_result[2]~q ),
	.datad(!\E_logic_result[2]~14_combout ),
	.datae(!\Add2~57_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[2]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[2]~15 .extended_lut = "off";
defparam \E_alu_result[2]~15 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_alu_result[2]~15 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_exception~0 (
	.dataa(!\Equal0~8_combout ),
	.datab(!\Equal0~9_combout ),
	.datac(!\Equal0~10_combout ),
	.datad(!\D_ctrl_exception~6_combout ),
	.datae(!\D_ctrl_exception~5_combout ),
	.dataf(!\D_ctrl_exception~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_exception~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_exception~0 .extended_lut = "off";
defparam \D_ctrl_exception~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \D_ctrl_exception~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_exception~3 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\D_iw[12]~q ),
	.datad(!\D_iw[11]~q ),
	.datae(!\D_iw[16]~q ),
	.dataf(!\D_iw[15]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_exception~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_exception~3 .extended_lut = "off";
defparam \D_ctrl_exception~3 .lut_mask = 64'hF7FFFFFFB3FFFFFF;
defparam \D_ctrl_exception~3 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_exception~2 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.datac(!\D_ctrl_exception~0_combout ),
	.datad(!\D_ctrl_exception~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_exception~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_exception~2 .extended_lut = "off";
defparam \D_ctrl_exception~2 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \D_ctrl_exception~2 .shared_arith = "off";

dffeas R_ctrl_exception(
	.clk(clk_clk),
	.d(\D_ctrl_exception~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_exception~q ),
	.prn(vcc));
defparam R_ctrl_exception.is_wysiwyg = "true";
defparam R_ctrl_exception.power_up = "low";

cyclonev_lcell_comb \D_ctrl_break~0 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[15]~q ),
	.datae(!\D_iw[16]~q ),
	.dataf(!\Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_break~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_break~0 .extended_lut = "off";
defparam \D_ctrl_break~0 .lut_mask = 64'hFBFFFFFFFFFFFFFF;
defparam \D_ctrl_break~0 .shared_arith = "off";

dffeas R_ctrl_break(
	.clk(clk_clk),
	.d(\D_ctrl_break~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_break~q ),
	.prn(vcc));
defparam R_ctrl_break.is_wysiwyg = "true";
defparam R_ctrl_break.power_up = "low";

cyclonev_lcell_comb \F_pc_sel_nxt.01~0 (
	.dataa(!\R_ctrl_exception~q ),
	.datab(!\R_ctrl_break~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_sel_nxt.01~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_sel_nxt.01~0 .extended_lut = "off";
defparam \F_pc_sel_nxt.01~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_pc_sel_nxt.01~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~12 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~12 .extended_lut = "off";
defparam \Equal0~12 .lut_mask = 64'hFFFFFFFFFFBFFFFF;
defparam \Equal0~12 .shared_arith = "off";

cyclonev_lcell_comb \Equal62~3 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~3 .extended_lut = "off";
defparam \Equal62~3 .lut_mask = 64'hFFFFFFFFFFFFFEFF;
defparam \Equal62~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~2 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~2 .extended_lut = "off";
defparam \Equal0~2 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \Equal0~2 .shared_arith = "off";

cyclonev_lcell_comb \E_invert_arith_src_msb~0 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal62~3_combout ),
	.datac(!\Equal0~1_combout ),
	.datad(!\Equal0~2_combout ),
	.datae(!\Equal62~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_invert_arith_src_msb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_invert_arith_src_msb~0 .extended_lut = "off";
defparam \E_invert_arith_src_msb~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \E_invert_arith_src_msb~0 .shared_arith = "off";

cyclonev_lcell_comb \E_invert_arith_src_msb~1 (
	.dataa(!\R_valid~q ),
	.datab(!\Equal0~6_combout ),
	.datac(!\Equal0~12_combout ),
	.datad(!\E_invert_arith_src_msb~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_invert_arith_src_msb~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_invert_arith_src_msb~1 .extended_lut = "off";
defparam \E_invert_arith_src_msb~1 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_invert_arith_src_msb~1 .shared_arith = "off";

dffeas E_invert_arith_src_msb(
	.clk(clk_clk),
	.d(\E_invert_arith_src_msb~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_invert_arith_src_msb~q ),
	.prn(vcc));
defparam E_invert_arith_src_msb.is_wysiwyg = "true";
defparam E_invert_arith_src_msb.power_up = "low";

cyclonev_lcell_comb \R_src2_hi[15]~13 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\R_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\R_src2_hi~1_combout ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[15]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[15]~13 .extended_lut = "off";
defparam \R_src2_hi[15]~13 .lut_mask = 64'hFF6FFFFFFF6FFFFF;
defparam \R_src2_hi[15]~13 .shared_arith = "off";

dffeas \E_src2[31] (
	.clk(clk_clk),
	.d(\R_src2_hi[15]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[31]~q ),
	.prn(vcc));
defparam \E_src2[31] .is_wysiwyg = "true";
defparam \E_src2[31] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[14]~14 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\R_ctrl_hi_imm16~q ),
	.datac(!\D_iw[20]~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[14]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[14]~14 .extended_lut = "off";
defparam \R_src2_hi[14]~14 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src2_hi[14]~14 .shared_arith = "off";

dffeas \E_src2[30] (
	.clk(clk_clk),
	.d(\R_src2_hi[14]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[30]~q ),
	.prn(vcc));
defparam \E_src2[30] .is_wysiwyg = "true";
defparam \E_src2[30] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[13]~16 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\R_ctrl_hi_imm16~q ),
	.datac(!\D_iw[19]~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[13]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[13]~16 .extended_lut = "off";
defparam \R_src2_hi[13]~16 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src2_hi[13]~16 .shared_arith = "off";

dffeas \E_src2[29] (
	.clk(clk_clk),
	.d(\R_src2_hi[13]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[29]~q ),
	.prn(vcc));
defparam \E_src2[29] .is_wysiwyg = "true";
defparam \E_src2[29] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[12]~15 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\R_ctrl_hi_imm16~q ),
	.datac(!\D_iw[18]~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[12]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[12]~15 .extended_lut = "off";
defparam \R_src2_hi[12]~15 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src2_hi[12]~15 .shared_arith = "off";

dffeas \E_src2[28] (
	.clk(clk_clk),
	.d(\R_src2_hi[12]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[28]~q ),
	.prn(vcc));
defparam \E_src2[28] .is_wysiwyg = "true";
defparam \E_src2[28] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[11]~3 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\R_ctrl_hi_imm16~q ),
	.datac(!\D_iw[17]~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[11]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[11]~3 .extended_lut = "off";
defparam \R_src2_hi[11]~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src2_hi[11]~3 .shared_arith = "off";

dffeas \E_src2[27] (
	.clk(clk_clk),
	.d(\R_src2_hi[11]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[27]~q ),
	.prn(vcc));
defparam \E_src2[27] .is_wysiwyg = "true";
defparam \E_src2[27] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[10]~12 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\R_src2_use_imm~q ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[10]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[10]~12 .extended_lut = "off";
defparam \R_src2_hi[10]~12 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src2_hi[10]~12 .shared_arith = "off";

dffeas \E_src2[26] (
	.clk(clk_clk),
	.d(\R_src2_hi[10]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[26]~q ),
	.prn(vcc));
defparam \E_src2[26] .is_wysiwyg = "true";
defparam \E_src2[26] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[9]~2 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\R_src2_use_imm~q ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[9]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[9]~2 .extended_lut = "off";
defparam \R_src2_hi[9]~2 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src2_hi[9]~2 .shared_arith = "off";

dffeas \E_src2[25] (
	.clk(clk_clk),
	.d(\R_src2_hi[9]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[25]~q ),
	.prn(vcc));
defparam \E_src2[25] .is_wysiwyg = "true";
defparam \E_src2[25] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[8]~9 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\R_src2_use_imm~q ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[8]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[8]~9 .extended_lut = "off";
defparam \R_src2_hi[8]~9 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src2_hi[8]~9 .shared_arith = "off";

dffeas \E_src2[24] (
	.clk(clk_clk),
	.d(\R_src2_hi[8]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[24]~q ),
	.prn(vcc));
defparam \E_src2[24] .is_wysiwyg = "true";
defparam \E_src2[24] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[7]~8 (
	.dataa(!\D_iw[13]~q ),
	.datab(!\R_src2_use_imm~q ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[7]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[7]~8 .extended_lut = "off";
defparam \R_src2_hi[7]~8 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src2_hi[7]~8 .shared_arith = "off";

dffeas \E_src2[23] (
	.clk(clk_clk),
	.d(\R_src2_hi[7]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[23]~q ),
	.prn(vcc));
defparam \E_src2[23] .is_wysiwyg = "true";
defparam \E_src2[23] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[6]~7 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\R_src2_use_imm~q ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[6]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[6]~7 .extended_lut = "off";
defparam \R_src2_hi[6]~7 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src2_hi[6]~7 .shared_arith = "off";

dffeas \E_src2[22] (
	.clk(clk_clk),
	.d(\R_src2_hi[6]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[22]~q ),
	.prn(vcc));
defparam \E_src2[22] .is_wysiwyg = "true";
defparam \E_src2[22] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[5]~6 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\R_src2_use_imm~q ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[5]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[5]~6 .extended_lut = "off";
defparam \R_src2_hi[5]~6 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src2_hi[5]~6 .shared_arith = "off";

dffeas \E_src2[21] (
	.clk(clk_clk),
	.d(\R_src2_hi[5]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[21]~q ),
	.prn(vcc));
defparam \E_src2[21] .is_wysiwyg = "true";
defparam \E_src2[21] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[4]~5 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\D_iw[10]~q ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[4]~5 .extended_lut = "off";
defparam \R_src2_hi[4]~5 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \R_src2_hi[4]~5 .shared_arith = "off";

dffeas \E_src2[20] (
	.clk(clk_clk),
	.d(\R_src2_hi[4]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[20]~q ),
	.prn(vcc));
defparam \E_src2[20] .is_wysiwyg = "true";
defparam \E_src2[20] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[3]~4 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\R_ctrl_hi_imm16~q ),
	.datac(!\D_iw[9]~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[3]~4 .extended_lut = "off";
defparam \R_src2_hi[3]~4 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src2_hi[3]~4 .shared_arith = "off";

dffeas \E_src2[19] (
	.clk(clk_clk),
	.d(\R_src2_hi[3]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[19]~q ),
	.prn(vcc));
defparam \E_src2[19] .is_wysiwyg = "true";
defparam \E_src2[19] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[2]~10 (
	.dataa(!\D_iw[8]~q ),
	.datab(!\R_src2_use_imm~q ),
	.datac(!\R_ctrl_hi_imm16~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[2]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[2]~10 .extended_lut = "off";
defparam \R_src2_hi[2]~10 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \R_src2_hi[2]~10 .shared_arith = "off";

dffeas \E_src2[18] (
	.clk(clk_clk),
	.d(\R_src2_hi[2]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[18]~q ),
	.prn(vcc));
defparam \E_src2[18] .is_wysiwyg = "true";
defparam \E_src2[18] .power_up = "low";

cyclonev_lcell_comb \R_src2_hi[1]~11 (
	.dataa(!\R_src2_use_imm~q ),
	.datab(!\R_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_iw[7]~q ),
	.datae(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\R_src2_hi[1]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \R_src2_hi[1]~11 .extended_lut = "off";
defparam \R_src2_hi[1]~11 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \R_src2_hi[1]~11 .shared_arith = "off";

dffeas \E_src2[17] (
	.clk(clk_clk),
	.d(\R_src2_hi[1]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[17]~q ),
	.prn(vcc));
defparam \E_src2[17] .is_wysiwyg = "true";
defparam \E_src2[17] .power_up = "low";

cyclonev_lcell_comb \Add2~65 (
	.dataa(gnd),
	.datab(!\E_alu_sub~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~65_sumout ),
	.cout(),
	.shareout());
defparam \Add2~65 .extended_lut = "off";
defparam \Add2~65 .lut_mask = 64'h0000000000003333;
defparam \Add2~65 .shared_arith = "off";

dffeas \R_compare_op[0] (
	.clk(clk_clk),
	.d(\D_logic_op_raw[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_compare_op[0]~q ),
	.prn(vcc));
defparam \R_compare_op[0] .is_wysiwyg = "true";
defparam \R_compare_op[0] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[25]~15 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[25]~q ),
	.datad(!\E_src1[25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[25]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[25]~15 .extended_lut = "off";
defparam \E_logic_result[25]~15 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[25]~15 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[27]~16 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[27]~q ),
	.datad(!\E_src1[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[27]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[27]~16 .extended_lut = "off";
defparam \E_logic_result[27]~16 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[27]~16 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~0 (
	.dataa(!\E_logic_result[25]~15_combout ),
	.datab(!\E_logic_result[27]~16_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~0 .extended_lut = "off";
defparam \Equal127~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Equal127~0 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[19]~17 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[19]~q ),
	.datad(!\E_src1[19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[19]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[19]~17 .extended_lut = "off";
defparam \E_logic_result[19]~17 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[19]~17 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[20]~18 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[20]~q ),
	.datad(!\E_src1[20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[20]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[20]~18 .extended_lut = "off";
defparam \E_logic_result[20]~18 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[20]~18 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[21]~19 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[21]~q ),
	.datad(!\E_src1[21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[21]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[21]~19 .extended_lut = "off";
defparam \E_logic_result[21]~19 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[21]~19 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[22]~20 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[22]~q ),
	.datad(!\E_src1[22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[22]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[22]~20 .extended_lut = "off";
defparam \E_logic_result[22]~20 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[22]~20 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[23]~21 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[23]~q ),
	.datad(!\E_src1[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[23]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[23]~21 .extended_lut = "off";
defparam \E_logic_result[23]~21 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[23]~21 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[24]~22 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[24]~q ),
	.datad(!\E_src1[24]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[24]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[24]~22 .extended_lut = "off";
defparam \E_logic_result[24]~22 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[24]~22 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~1 (
	.dataa(!\E_logic_result[19]~17_combout ),
	.datab(!\E_logic_result[20]~18_combout ),
	.datac(!\E_logic_result[21]~19_combout ),
	.datad(!\E_logic_result[22]~20_combout ),
	.datae(!\E_logic_result[23]~21_combout ),
	.dataf(!\E_logic_result[24]~22_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~1 .extended_lut = "off";
defparam \Equal127~1 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal127~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~2 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[14]~q ),
	.datad(!\E_src2[14]~q ),
	.datae(!\E_src1[15]~q ),
	.dataf(!\E_src2[15]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~2 .extended_lut = "off";
defparam \Equal127~2 .lut_mask = 64'h6996966996696996;
defparam \Equal127~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~3 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[12]~q ),
	.datad(!\E_src2[12]~q ),
	.datae(!\E_src1[13]~q ),
	.dataf(!\E_src2[13]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~3 .extended_lut = "off";
defparam \Equal127~3 .lut_mask = 64'h6996966996696996;
defparam \Equal127~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~4 (
	.dataa(!\E_src1[4]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\R_logic_op[1]~q ),
	.datad(!\R_logic_op[0]~q ),
	.datae(!\E_src2[5]~q ),
	.dataf(!\E_src1[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~4 .extended_lut = "off";
defparam \Equal127~4 .lut_mask = 64'h6996966996696996;
defparam \Equal127~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~5 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[7]~q ),
	.datad(!\E_src1[7]~q ),
	.datae(!\E_src2[6]~q ),
	.dataf(!\E_src1[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~5 .extended_lut = "off";
defparam \Equal127~5 .lut_mask = 64'h6996966996696996;
defparam \Equal127~5 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~6 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src1[11]~q ),
	.datad(!\E_src2[11]~q ),
	.datae(!\E_src2[10]~q ),
	.dataf(!\E_src1[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~6 .extended_lut = "off";
defparam \Equal127~6 .lut_mask = 64'h6996966996696996;
defparam \Equal127~6 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~7 (
	.dataa(!\E_logic_result[9]~3_combout ),
	.datab(!\E_logic_result[8]~4_combout ),
	.datac(!\Equal127~3_combout ),
	.datad(!\Equal127~4_combout ),
	.datae(!\Equal127~5_combout ),
	.dataf(!\Equal127~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~7 .extended_lut = "off";
defparam \Equal127~7 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \Equal127~7 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~8 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[18]~q ),
	.datad(!\E_src1[18]~q ),
	.datae(!\E_src2[17]~q ),
	.dataf(!\E_src1[17]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~8 .extended_lut = "off";
defparam \Equal127~8 .lut_mask = 64'h6996966996696996;
defparam \Equal127~8 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~9 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[1]~q ),
	.datad(!\E_src1[1]~q ),
	.datae(!\E_src2[26]~q ),
	.dataf(!\E_src1[26]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~9 .extended_lut = "off";
defparam \Equal127~9 .lut_mask = 64'h6996966996696996;
defparam \Equal127~9 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~10 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[31]~q ),
	.datad(!\E_src1[31]~q ),
	.datae(!\E_src2[30]~q ),
	.dataf(!\E_src1[30]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~10 .extended_lut = "off";
defparam \Equal127~10 .lut_mask = 64'h6996966996696996;
defparam \Equal127~10 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[0]~23 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_src1[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[0]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[0]~23 .extended_lut = "off";
defparam \E_logic_result[0]~23 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[0]~23 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[28]~24 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[28]~q ),
	.datad(!\E_src1[28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[28]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[28]~24 .extended_lut = "off";
defparam \E_logic_result[28]~24 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[28]~24 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[29]~25 (
	.dataa(!\R_logic_op[1]~q ),
	.datab(!\R_logic_op[0]~q ),
	.datac(!\E_src2[29]~q ),
	.datad(!\E_src1[29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[29]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[29]~25 .extended_lut = "off";
defparam \E_logic_result[29]~25 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[29]~25 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~11 (
	.dataa(!\E_logic_result[16]~12_combout ),
	.datab(!\E_logic_result[3]~13_combout ),
	.datac(!\E_logic_result[2]~14_combout ),
	.datad(!\E_logic_result[0]~23_combout ),
	.datae(!\E_logic_result[28]~24_combout ),
	.dataf(!\E_logic_result[29]~25_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~11 .extended_lut = "off";
defparam \Equal127~11 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal127~11 .shared_arith = "off";

cyclonev_lcell_comb \Equal127~12 (
	.dataa(!\Equal127~2_combout ),
	.datab(!\Equal127~7_combout ),
	.datac(!\Equal127~8_combout ),
	.datad(!\Equal127~9_combout ),
	.datae(!\Equal127~10_combout ),
	.dataf(!\Equal127~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal127~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal127~12 .extended_lut = "off";
defparam \Equal127~12 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \Equal127~12 .shared_arith = "off";

dffeas \R_compare_op[1] (
	.clk(clk_clk),
	.d(\D_logic_op_raw[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_compare_op[1]~q ),
	.prn(vcc));
defparam \R_compare_op[1] .is_wysiwyg = "true";
defparam \R_compare_op[1] .power_up = "low";

cyclonev_lcell_comb \E_cmp_result~0 (
	.dataa(!\Add2~65_sumout ),
	.datab(!\R_compare_op[0]~q ),
	.datac(!\Equal127~0_combout ),
	.datad(!\Equal127~1_combout ),
	.datae(!\Equal127~12_combout ),
	.dataf(!\R_compare_op[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_cmp_result~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_cmp_result~0 .extended_lut = "off";
defparam \E_cmp_result~0 .lut_mask = 64'h6996966996696996;
defparam \E_cmp_result~0 .shared_arith = "off";

dffeas W_cmp_result(
	.clk(clk_clk),
	.d(\E_cmp_result~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_cmp_result~q ),
	.prn(vcc));
defparam W_cmp_result.is_wysiwyg = "true";
defparam W_cmp_result.power_up = "low";

cyclonev_lcell_comb \Equal62~12 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal62~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal62~12 .extended_lut = "off";
defparam \Equal62~12 .lut_mask = 64'hFFFFFFFFDFFFFFFF;
defparam \Equal62~12 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_uncond_cti_non_br~0 (
	.dataa(!\Equal62~12_combout ),
	.datab(!\Equal62~13_combout ),
	.datac(!\Equal62~14_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_uncond_cti_non_br~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_uncond_cti_non_br~0 .extended_lut = "off";
defparam \D_ctrl_uncond_cti_non_br~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \D_ctrl_uncond_cti_non_br~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_uncond_cti_non_br~1 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal62~15_combout ),
	.datac(!\Equal62~16_combout ),
	.datad(!\D_ctrl_uncond_cti_non_br~0_combout ),
	.datae(!\D_ctrl_jmp_direct~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_uncond_cti_non_br~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_uncond_cti_non_br~1 .extended_lut = "off";
defparam \D_ctrl_uncond_cti_non_br~1 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \D_ctrl_uncond_cti_non_br~1 .shared_arith = "off";

dffeas R_ctrl_uncond_cti_non_br(
	.clk(clk_clk),
	.d(\D_ctrl_uncond_cti_non_br~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_uncond_cti_non_br~q ),
	.prn(vcc));
defparam R_ctrl_uncond_cti_non_br.is_wysiwyg = "true";
defparam R_ctrl_uncond_cti_non_br.power_up = "low";

cyclonev_lcell_comb \Equal0~3 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~3 .extended_lut = "off";
defparam \Equal0~3 .lut_mask = 64'hFFFFFFFFFFFFFFBF;
defparam \Equal0~3 .shared_arith = "off";

dffeas R_ctrl_br_uncond(
	.clk(clk_clk),
	.d(\Equal0~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br_uncond~q ),
	.prn(vcc));
defparam R_ctrl_br_uncond.is_wysiwyg = "true";
defparam R_ctrl_br_uncond.power_up = "low";

cyclonev_lcell_comb \F_pc_sel_nxt~0 (
	.dataa(!\W_cmp_result~q ),
	.datab(!\R_ctrl_br~q ),
	.datac(!\R_ctrl_uncond_cti_non_br~q ),
	.datad(!\R_ctrl_br_uncond~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_sel_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_sel_nxt~0 .extended_lut = "off";
defparam \F_pc_sel_nxt~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \F_pc_sel_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_sel_nxt.10~0 (
	.dataa(!\R_ctrl_exception~q ),
	.datab(!\R_ctrl_break~q ),
	.datac(!\F_pc_sel_nxt~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_sel_nxt.10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_sel_nxt.10~0 .extended_lut = "off";
defparam \F_pc_sel_nxt.10~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \F_pc_sel_nxt.10~0 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[9]~0 (
	.dataa(!\Add2~5_sumout ),
	.datab(!\Add0~5_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[9]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[9]~0 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[9]~0 .lut_mask = 64'h5F3F5F3F5F3F5F3F;
defparam \F_pc_no_crst_nxt[9]~0 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[10]~1 (
	.dataa(!\Add2~33_sumout ),
	.datab(!\Add0~33_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[10]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[10]~1 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[10]~1 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[10]~1 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[11]~2 (
	.dataa(!\Add2~37_sumout ),
	.datab(!\Add0~37_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[11]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[11]~2 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[11]~2 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[11]~2 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[12]~3 (
	.dataa(!\Add2~41_sumout ),
	.datab(!\Add0~41_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[12]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[12]~3 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[12]~3 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[12]~3 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[14]~5 (
	.dataa(!\Add2~49_sumout ),
	.datab(!\Add0~49_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[14]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[14]~5 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[14]~5 .lut_mask = 64'h5F3F5F3F5F3F5F3F;
defparam \F_pc_no_crst_nxt[14]~5 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[2]~6 (
	.dataa(!\Add2~1_sumout ),
	.datab(!\Add0~1_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[2]~6 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[2]~6 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[8]~7 (
	.dataa(!\Add2~9_sumout ),
	.datab(!\Add0~9_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[8]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[8]~7 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[8]~7 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[8]~7 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[7]~8 (
	.dataa(!\Add2~13_sumout ),
	.datab(!\Add0~13_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[7]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[7]~8 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[7]~8 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[7]~8 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[6]~9 (
	.dataa(!\Add2~17_sumout ),
	.datab(!\Add0~17_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[6]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[6]~9 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[6]~9 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[6]~9 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[5]~10 (
	.dataa(!\Add2~21_sumout ),
	.datab(!\Add0~21_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[5]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[5]~10 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[5]~10 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[5]~10 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[4]~11 (
	.dataa(!\Add2~25_sumout ),
	.datab(!\Add0~25_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[4]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[4]~11 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[4]~11 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[4]~11 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt~12 (
	.dataa(!\Add2~29_sumout ),
	.datab(!\Add0~29_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt~12 .extended_lut = "off";
defparam \F_pc_no_crst_nxt~12 .lut_mask = 64'h5F3F5F3F5F3F5F3F;
defparam \F_pc_no_crst_nxt~12 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[1]~13 (
	.dataa(!\Add2~53_sumout ),
	.datab(!\Add0~53_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[1]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[1]~13 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[1]~13 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[1]~13 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[0]~14 (
	.dataa(!\Add2~57_sumout ),
	.datab(!\Add0~57_sumout ),
	.datac(!\F_pc_sel_nxt.01~0_combout ),
	.datad(!\F_pc_sel_nxt.10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[0]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[0]~14 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[0]~14 .lut_mask = 64'hF377F377F377F377;
defparam \F_pc_no_crst_nxt[0]~14 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_mem8~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_mem8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_mem8~0 .extended_lut = "off";
defparam \D_ctrl_mem8~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \D_ctrl_mem8~0 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[23]~0 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_ctrl_mem16~0_combout ),
	.datac(!\D_ctrl_mem8~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[23]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[23]~0 .extended_lut = "off";
defparam \E_st_data[23]~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \E_st_data[23]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_mem8~1 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_ctrl_mem8~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_mem8~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_mem8~1 .extended_lut = "off";
defparam \D_ctrl_mem8~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \D_ctrl_mem8~1 .shared_arith = "off";

cyclonev_lcell_comb E_st_stall(
	.dataa(!d_write1),
	.datab(!\d_write_nxt~0_combout ),
	.datac(!av_waitrequest1),
	.datad(!read_latency_shift_reg),
	.datae(!WideOr0),
	.dataf(!av_waitrequest),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_stall~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_st_stall.extended_lut = "off";
defparam E_st_stall.lut_mask = 64'hFF7FFFFFFFFFFFFF;
defparam E_st_stall.shared_arith = "off";

cyclonev_lcell_comb d_read_nxt(
	.dataa(!d_read1),
	.datab(!\E_new_inst~q ),
	.datac(!src0_valid),
	.datad(!WideOr1),
	.datae(!\R_ctrl_ld~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_read_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam d_read_nxt.extended_lut = "off";
defparam d_read_nxt.lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam d_read_nxt.shared_arith = "off";

cyclonev_lcell_comb \i_read_nxt~0 (
	.dataa(!\W_valid~q ),
	.datab(!i_read1),
	.datac(!src1_valid1),
	.datad(!src1_valid2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\i_read_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \i_read_nxt~0 .extended_lut = "off";
defparam \i_read_nxt~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \i_read_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_no_crst_nxt[13]~4 (
	.dataa(!\Add2~45_sumout ),
	.datab(!\Add0~45_sumout ),
	.datac(!\R_ctrl_exception~q ),
	.datad(!\R_ctrl_break~q ),
	.datae(!\F_pc_sel_nxt~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_no_crst_nxt[13]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_no_crst_nxt[13]~4 .extended_lut = "off";
defparam \F_pc_no_crst_nxt[13]~4 .lut_mask = 64'hFAFFFCFFFAFFFCFF;
defparam \F_pc_no_crst_nxt[13]~4 .shared_arith = "off";

cyclonev_lcell_comb \hbreak_enabled~0 (
	.dataa(!\Equal0~0_combout ),
	.datab(!hbreak_enabled1),
	.datac(!\Equal62~16_combout ),
	.datad(!\R_ctrl_break~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hbreak_enabled~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hbreak_enabled~0 .extended_lut = "off";
defparam \hbreak_enabled~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \hbreak_enabled~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_mem16~1 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_ctrl_mem16~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_mem16~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_mem16~1 .extended_lut = "off";
defparam \D_ctrl_mem16~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \D_ctrl_mem16~1 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en~0 (
	.dataa(!\Add2~61_sumout ),
	.datab(!\D_ctrl_mem16~1_combout ),
	.datac(!\Add2~69_sumout ),
	.datad(!\D_ctrl_mem8~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en~0 .extended_lut = "off";
defparam \E_mem_byte_en~0 .lut_mask = 64'hFBFEFBFEFBFEFBFE;
defparam \E_mem_byte_en~0 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en[2]~1 (
	.dataa(!\Add2~61_sumout ),
	.datab(!\D_ctrl_mem16~1_combout ),
	.datac(!\Add2~69_sumout ),
	.datad(!\D_ctrl_mem8~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en[2]~1 .extended_lut = "off";
defparam \E_mem_byte_en[2]~1 .lut_mask = 64'hF7FDF7FDF7FDF7FD;
defparam \E_mem_byte_en[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[24]~1 (
	.dataa(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datab(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datac(!\D_ctrl_mem16~1_combout ),
	.datad(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.datae(!\D_ctrl_mem8~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[24]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[24]~1 .extended_lut = "off";
defparam \E_st_data[24]~1 .lut_mask = 64'h7FFFF7FF7FFFF7FF;
defparam \E_st_data[24]~1 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en[3]~2 (
	.dataa(!\Add2~61_sumout ),
	.datab(!\D_ctrl_mem16~1_combout ),
	.datac(!\Add2~69_sumout ),
	.datad(!\D_ctrl_mem8~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en[3]~2 .extended_lut = "off";
defparam \E_mem_byte_en[3]~2 .lut_mask = 64'h7FDF7FDF7FDF7FDF;
defparam \E_mem_byte_en[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[25]~2 (
	.dataa(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datab(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datac(!\D_ctrl_mem16~1_combout ),
	.datad(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.datae(!\D_ctrl_mem8~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[25]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[25]~2 .extended_lut = "off";
defparam \E_st_data[25]~2 .lut_mask = 64'h7FFFF7FF7FFFF7FF;
defparam \E_st_data[25]~2 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[26]~3 (
	.dataa(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datab(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datac(!\D_ctrl_mem16~1_combout ),
	.datad(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.datae(!\D_ctrl_mem8~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[26]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[26]~3 .extended_lut = "off";
defparam \E_st_data[26]~3 .lut_mask = 64'h7FFFF7FF7FFFF7FF;
defparam \E_st_data[26]~3 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en[1]~3 (
	.dataa(!\Add2~61_sumout ),
	.datab(!\D_ctrl_mem16~1_combout ),
	.datac(!\Add2~69_sumout ),
	.datad(!\D_ctrl_mem8~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en[1]~3 .extended_lut = "off";
defparam \E_mem_byte_en[1]~3 .lut_mask = 64'hBFEFBFEFBFEFBFEF;
defparam \E_mem_byte_en[1]~3 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[27]~4 (
	.dataa(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datab(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datac(!\D_ctrl_mem16~1_combout ),
	.datad(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.datae(!\D_ctrl_mem8~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[27]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[27]~4 .extended_lut = "off";
defparam \E_st_data[27]~4 .lut_mask = 64'h7FFFF7FF7FFFF7FF;
defparam \E_st_data[27]~4 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[28]~5 (
	.dataa(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datab(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datac(!\D_ctrl_mem16~1_combout ),
	.datad(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.datae(!\D_ctrl_mem8~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[28]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[28]~5 .extended_lut = "off";
defparam \E_st_data[28]~5 .lut_mask = 64'h7FFFF7FF7FFFF7FF;
defparam \E_st_data[28]~5 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[29]~6 (
	.dataa(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.datab(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datac(!\D_ctrl_mem16~1_combout ),
	.datad(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.datae(!\D_ctrl_mem8~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[29]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[29]~6 .extended_lut = "off";
defparam \E_st_data[29]~6 .lut_mask = 64'h7FFFF7FF7FFFF7FF;
defparam \E_st_data[29]~6 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[30]~7 (
	.dataa(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.datab(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datac(!\D_ctrl_mem16~1_combout ),
	.datad(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.datae(!\D_ctrl_mem8~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[30]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[30]~7 .extended_lut = "off";
defparam \E_st_data[30]~7 .lut_mask = 64'h7FFFF7FF7FFFF7FF;
defparam \E_st_data[30]~7 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[31]~8 (
	.dataa(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.datab(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datac(!\D_ctrl_mem16~1_combout ),
	.datad(!\niosLab2_nios2_gen2_0_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.datae(!\D_ctrl_mem8~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[31]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[31]~8 .extended_lut = "off";
defparam \E_st_data[31]~8 .lut_mask = 64'h7FFFF7FF7FFFF7FF;
defparam \E_st_data[31]~8 .shared_arith = "off";

endmodule

module niosLab2_niosLab2_nios2_gen2_0_cpu_nios2_oci (
	readdata_0,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_11,
	readdata_12,
	readdata_13,
	readdata_14,
	readdata_15,
	readdata_16,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_8,
	readdata_10,
	readdata_17,
	readdata_9,
	readdata_18,
	readdata_19,
	readdata_20,
	readdata_21,
	readdata_6,
	readdata_7,
	readdata_27,
	readdata_28,
	readdata_29,
	readdata_30,
	readdata_31,
	sr_0,
	ir_out_0,
	ir_out_1,
	r_sync_rst,
	always2,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	src1_valid,
	src_valid,
	mem,
	hbreak_enabled,
	jtag_break,
	address_nxt,
	r_early_rst,
	oci_single_step_mode,
	writedata_nxt,
	debugaccess_nxt,
	byteenable_nxt,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	readdata_0;
output 	readdata_22;
output 	readdata_23;
output 	readdata_24;
output 	readdata_25;
output 	readdata_26;
output 	readdata_11;
output 	readdata_12;
output 	readdata_13;
output 	readdata_14;
output 	readdata_15;
output 	readdata_16;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_8;
output 	readdata_10;
output 	readdata_17;
output 	readdata_9;
output 	readdata_18;
output 	readdata_19;
output 	readdata_20;
output 	readdata_21;
output 	readdata_6;
output 	readdata_7;
output 	readdata_27;
output 	readdata_28;
output 	readdata_29;
output 	readdata_30;
output 	readdata_31;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	r_sync_rst;
input 	always2;
input 	saved_grant_0;
output 	waitrequest;
input 	mem_used_1;
input 	src1_valid;
input 	src_valid;
input 	mem;
input 	hbreak_enabled;
output 	jtag_break;
input 	[8:0] address_nxt;
input 	r_early_rst;
output 	oci_single_step_mode;
input 	[31:0] writedata_nxt;
input 	debugaccess_nxt;
input 	[3:0] byteenable_nxt;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[0]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[1]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[1]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[2]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[2]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[3]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[3]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[16]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[16]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[24]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[24]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[4]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[25]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[25]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[27]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[27]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[26]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[26]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[22]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[20]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[20]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[19]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[19]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[23]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[11]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[13]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[14]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[10]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[17]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[9]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[21]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[6]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[17]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[7]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[5]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[28]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[28]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[29]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[30]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[30]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[31]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[31]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[21]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[18]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[6]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[22]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[15]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[23]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[7]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[13]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[14]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[10]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[12]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[11]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[8]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[9]~q ;
wire \read~0_combout ;
wire \write~0_combout ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[0]~q ;
wire \write~q ;
wire \read~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug|monitor_ready~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[0]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[36]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[37]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|ir[1]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|ir[0]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|enable_action_strobe~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[35]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[3]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[34]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[17]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[25]~q ;
wire \writedata[0]~q ;
wire \address[3]~q ;
wire \address[7]~q ;
wire \address[6]~q ;
wire \address[5]~q ;
wire \address[4]~q ;
wire \address[2]~q ;
wire \address[1]~q ;
wire \debugaccess~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[1]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[4]~q ;
wire \byteenable[0]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[26]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[28]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[27]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[21]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[20]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[2]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[5]~q ;
wire \writedata[1]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[29]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[30]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[31]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[32]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[33]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|Equal0~2_combout ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug|monitor_error~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[19]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[18]~q ;
wire \writedata[3]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug|monitor_go~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[4]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[6]~q ;
wire \writedata[2]~q ;
wire \writedata[22]~q ;
wire \byteenable[2]~q ;
wire \writedata[23]~q ;
wire \writedata[24]~q ;
wire \byteenable[3]~q ;
wire \writedata[25]~q ;
wire \writedata[26]~q ;
wire \writedata[11]~q ;
wire \byteenable[1]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[12]~q ;
wire \writedata[12]~q ;
wire \writedata[13]~q ;
wire \writedata[14]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[15]~q ;
wire \writedata[15]~q ;
wire \writedata[16]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[23]~q ;
wire \writedata[4]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[5]~q ;
wire \writedata[5]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[8]~q ;
wire \writedata[8]~q ;
wire \writedata[10]~q ;
wire \writedata[17]~q ;
wire \writedata[9]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[18]~q ;
wire \writedata[18]~q ;
wire \writedata[19]~q ;
wire \writedata[20]~q ;
wire \writedata[21]~q ;
wire \writedata[6]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[16]~q ;
wire \writedata[7]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[24]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[7]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[29]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug|resetlatch~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[22]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[14]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[15]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[8]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[11]~q ;
wire \writedata[27]~q ;
wire \writedata[28]~q ;
wire \writedata[29]~q ;
wire \writedata[30]~q ;
wire \writedata[31]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[13]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[12]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[9]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[10]~q ;
wire \address[0]~q ;
wire \readdata~0_combout ;
wire \address[8]~q ;
wire \readdata~1_combout ;
wire \readdata~2_combout ;
wire \readdata~3_combout ;


niosLab2_niosLab2_nios2_gen2_0_cpu_nios2_oci_break the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break(
	.break_readreg_0(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[0]~q ),
	.break_readreg_1(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[1]~q ),
	.break_readreg_2(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[2]~q ),
	.break_readreg_3(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[3]~q ),
	.break_readreg_16(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[16]~q ),
	.break_readreg_24(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[24]~q ),
	.break_readreg_4(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[4]~q ),
	.break_readreg_25(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[25]~q ),
	.break_readreg_27(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[27]~q ),
	.break_readreg_26(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[26]~q ),
	.break_readreg_20(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[20]~q ),
	.break_readreg_19(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[19]~q ),
	.break_readreg_17(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[17]~q ),
	.break_readreg_5(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[5]~q ),
	.break_readreg_28(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[28]~q ),
	.break_readreg_29(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[29]~q ),
	.break_readreg_30(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[30]~q ),
	.break_readreg_31(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[31]~q ),
	.break_readreg_21(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[21]~q ),
	.break_readreg_18(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_6(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[6]~q ),
	.break_readreg_22(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[22]~q ),
	.break_readreg_15(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_23(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[23]~q ),
	.break_readreg_7(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_13(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_14(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_10(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_12(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_11(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[11]~q ),
	.break_readreg_8(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[8]~q ),
	.break_readreg_9(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[9]~q ),
	.jdo_0(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[0]~q ),
	.jdo_36(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[36]~q ),
	.jdo_37(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[37]~q ),
	.ir_1(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|ir[1]~q ),
	.ir_0(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|ir[0]~q ),
	.enable_action_strobe(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|enable_action_strobe~q ),
	.jdo_3(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[3]~q ),
	.jdo_17(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[17]~q ),
	.jdo_25(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_1(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[1]~q ),
	.jdo_4(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_28(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_21(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[20]~q ),
	.jdo_2(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[2]~q ),
	.jdo_5(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[5]~q ),
	.jdo_29(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_30(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_31(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_19(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[18]~q ),
	.jdo_6(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[6]~q ),
	.jdo_23(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[23]~q ),
	.jdo_16(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[16]~q ),
	.jdo_24(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[24]~q ),
	.jdo_7(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[7]~q ),
	.jdo_22(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_14(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_8(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_11(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_13(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_9(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[9]~q ),
	.jdo_10(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[10]~q ),
	.clk_clk(clk_clk));

niosLab2_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug the_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug(
	.r_sync_rst(r_sync_rst),
	.monitor_ready1(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug|monitor_ready~q ),
	.jtag_break1(jtag_break),
	.jdo_34(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[34]~q ),
	.take_action_ocimem_a(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ),
	.take_action_ocimem_a1(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.jdo_25(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[25]~q ),
	.writedata_0(\writedata[0]~q ),
	.take_action_ocireg(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.jdo_21(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[20]~q ),
	.writedata_1(\writedata[1]~q ),
	.monitor_error1(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug|monitor_error~q ),
	.jdo_19(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[18]~q ),
	.monitor_go1(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug|monitor_go~q ),
	.jdo_23(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[23]~q ),
	.jdo_24(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[24]~q ),
	.resetlatch1(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug|resetlatch~q ),
	.state_1(state_1),
	.clk_clk(clk_clk));

niosLab2_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper(
	.break_readreg_0(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[0]~q ),
	.break_readreg_1(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[1]~q ),
	.MonDReg_1(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[1]~q ),
	.break_readreg_2(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[2]~q ),
	.MonDReg_2(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[2]~q ),
	.break_readreg_3(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[3]~q ),
	.MonDReg_3(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[3]~q ),
	.break_readreg_16(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[16]~q ),
	.MonDReg_16(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[16]~q ),
	.break_readreg_24(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[24]~q ),
	.MonDReg_24(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[24]~q ),
	.break_readreg_4(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[4]~q ),
	.break_readreg_25(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[25]~q ),
	.MonDReg_25(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[25]~q ),
	.break_readreg_27(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[27]~q ),
	.MonDReg_27(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[27]~q ),
	.break_readreg_26(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[26]~q ),
	.MonDReg_26(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[26]~q ),
	.MonDReg_22(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[22]~q ),
	.break_readreg_20(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[20]~q ),
	.MonDReg_20(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[20]~q ),
	.break_readreg_19(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[19]~q ),
	.MonDReg_19(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[19]~q ),
	.MonDReg_23(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[23]~q ),
	.MonDReg_11(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[11]~q ),
	.MonDReg_13(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[13]~q ),
	.MonDReg_14(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[14]~q ),
	.MonDReg_10(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[10]~q ),
	.MonDReg_17(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[17]~q ),
	.MonDReg_9(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[9]~q ),
	.MonDReg_21(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[21]~q ),
	.MonDReg_6(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[6]~q ),
	.break_readreg_17(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[17]~q ),
	.MonDReg_7(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[7]~q ),
	.break_readreg_5(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[5]~q ),
	.break_readreg_28(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[28]~q ),
	.MonDReg_28(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[28]~q ),
	.break_readreg_29(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[29]~q ),
	.MonDReg_30(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[30]~q ),
	.break_readreg_30(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[30]~q ),
	.break_readreg_31(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[31]~q ),
	.MonDReg_31(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[31]~q ),
	.break_readreg_21(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[21]~q ),
	.break_readreg_18(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_6(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[6]~q ),
	.break_readreg_22(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[22]~q ),
	.break_readreg_15(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_23(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[23]~q ),
	.break_readreg_7(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_13(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_14(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_10(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_12(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_11(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[11]~q ),
	.break_readreg_8(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[8]~q ),
	.break_readreg_9(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_break|break_readreg[9]~q ),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.MonDReg_0(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[0]~q ),
	.monitor_ready(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug|monitor_ready~q ),
	.jdo_0(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[0]~q ),
	.jdo_36(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[36]~q ),
	.jdo_37(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[37]~q ),
	.ir_1(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|ir[1]~q ),
	.ir_0(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|ir[0]~q ),
	.enable_action_strobe(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|enable_action_strobe~q ),
	.jdo_35(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[35]~q ),
	.take_action_ocimem_b(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ),
	.jdo_3(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[3]~q ),
	.hbreak_enabled(hbreak_enabled),
	.take_action_ocimem_a(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.jdo_34(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[34]~q ),
	.jdo_17(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[17]~q ),
	.take_action_ocimem_a1(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ),
	.take_action_ocimem_a2(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.jdo_25(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_1(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[1]~q ),
	.jdo_4(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_26(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_28(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_21(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[20]~q ),
	.jdo_2(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[2]~q ),
	.jdo_5(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[5]~q ),
	.jdo_29(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_30(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_31(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_32(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[32]~q ),
	.jdo_33(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[33]~q ),
	.monitor_error(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug|monitor_error~q ),
	.jdo_19(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[18]~q ),
	.MonDReg_4(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[4]~q ),
	.jdo_6(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[6]~q ),
	.MonDReg_12(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[12]~q ),
	.MonDReg_15(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[15]~q ),
	.jdo_23(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[23]~q ),
	.MonDReg_5(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[5]~q ),
	.MonDReg_8(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[8]~q ),
	.MonDReg_18(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[18]~q ),
	.jdo_16(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[16]~q ),
	.jdo_24(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[24]~q ),
	.jdo_7(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[7]~q ),
	.MonDReg_29(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[29]~q ),
	.resetlatch(\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug|resetlatch~q ),
	.jdo_22(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_14(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_8(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_11(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_13(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_9(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[9]~q ),
	.jdo_10(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[10]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

niosLab2_niosLab2_nios2_gen2_0_cpu_nios2_ocimem the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem(
	.MonDReg_1(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[1]~q ),
	.q_a_0(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.MonDReg_2(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[2]~q ),
	.q_a_1(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.MonDReg_3(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[3]~q ),
	.q_a_2(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_22(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_23(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_24(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_25(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_26(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_11(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_12(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_13(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_14(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_15(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_16(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_3(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_4(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_5(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_8(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_10(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_17(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_9(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_18(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_19(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_20(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_21(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_6(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.MonDReg_16(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[16]~q ),
	.q_a_7(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.MonDReg_24(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[24]~q ),
	.MonDReg_25(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[25]~q ),
	.MonDReg_27(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[27]~q ),
	.MonDReg_26(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[26]~q ),
	.MonDReg_22(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[22]~q ),
	.MonDReg_20(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[20]~q ),
	.MonDReg_19(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[19]~q ),
	.MonDReg_23(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[23]~q ),
	.MonDReg_11(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[11]~q ),
	.MonDReg_13(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[13]~q ),
	.MonDReg_14(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[14]~q ),
	.q_a_27(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_28(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_29(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_30(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_31(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.MonDReg_10(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[10]~q ),
	.MonDReg_17(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[17]~q ),
	.MonDReg_9(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[9]~q ),
	.MonDReg_21(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[21]~q ),
	.MonDReg_6(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[6]~q ),
	.MonDReg_7(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[7]~q ),
	.MonDReg_28(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[28]~q ),
	.MonDReg_30(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[30]~q ),
	.MonDReg_31(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[31]~q ),
	.waitrequest1(waitrequest),
	.MonDReg_0(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[0]~q ),
	.write(\write~q ),
	.address_8(\address[8]~q ),
	.read(\read~q ),
	.ir_1(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|ir[1]~q ),
	.ir_0(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|ir[0]~q ),
	.enable_action_strobe(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|enable_action_strobe~q ),
	.jdo_35(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[35]~q ),
	.take_action_ocimem_b(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ),
	.jdo_3(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[3]~q ),
	.take_action_ocimem_a(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.jdo_34(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[34]~q ),
	.jdo_17(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[17]~q ),
	.take_action_ocimem_a1(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ),
	.take_action_ocimem_a2(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.jdo_25(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[25]~q ),
	.writedata_0(\writedata[0]~q ),
	.address_0(\address[0]~q ),
	.address_3(\address[3]~q ),
	.address_7(\address[7]~q ),
	.address_6(\address[6]~q ),
	.address_5(\address[5]~q ),
	.address_4(\address[4]~q ),
	.address_2(\address[2]~q ),
	.address_1(\address[1]~q ),
	.debugaccess(\debugaccess~q ),
	.jdo_4(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[4]~q ),
	.r_early_rst(r_early_rst),
	.byteenable_0(\byteenable[0]~q ),
	.jdo_26(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[26]~q ),
	.jdo_28(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_21(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[20]~q ),
	.jdo_5(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[5]~q ),
	.writedata_1(\writedata[1]~q ),
	.jdo_29(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_30(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_31(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_32(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[32]~q ),
	.jdo_33(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[33]~q ),
	.jdo_19(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[18]~q ),
	.writedata_3(\writedata[3]~q ),
	.MonDReg_4(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[4]~q ),
	.jdo_6(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[6]~q ),
	.writedata_2(\writedata[2]~q ),
	.writedata_22(\writedata[22]~q ),
	.byteenable_2(\byteenable[2]~q ),
	.writedata_23(\writedata[23]~q ),
	.writedata_24(\writedata[24]~q ),
	.byteenable_3(\byteenable[3]~q ),
	.writedata_25(\writedata[25]~q ),
	.writedata_26(\writedata[26]~q ),
	.writedata_11(\writedata[11]~q ),
	.byteenable_1(\byteenable[1]~q ),
	.MonDReg_12(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[12]~q ),
	.writedata_12(\writedata[12]~q ),
	.writedata_13(\writedata[13]~q ),
	.writedata_14(\writedata[14]~q ),
	.MonDReg_15(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[15]~q ),
	.writedata_15(\writedata[15]~q ),
	.writedata_16(\writedata[16]~q ),
	.jdo_23(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[23]~q ),
	.writedata_4(\writedata[4]~q ),
	.MonDReg_5(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[5]~q ),
	.writedata_5(\writedata[5]~q ),
	.MonDReg_8(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[8]~q ),
	.writedata_8(\writedata[8]~q ),
	.writedata_10(\writedata[10]~q ),
	.writedata_17(\writedata[17]~q ),
	.writedata_9(\writedata[9]~q ),
	.MonDReg_18(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[18]~q ),
	.writedata_18(\writedata[18]~q ),
	.writedata_19(\writedata[19]~q ),
	.writedata_20(\writedata[20]~q ),
	.writedata_21(\writedata[21]~q ),
	.writedata_6(\writedata[6]~q ),
	.jdo_16(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[16]~q ),
	.writedata_7(\writedata[7]~q ),
	.jdo_24(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[24]~q ),
	.jdo_7(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[7]~q ),
	.MonDReg_29(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|MonDReg[29]~q ),
	.jdo_22(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_14(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_8(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_11(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[11]~q ),
	.writedata_27(\writedata[27]~q ),
	.writedata_28(\writedata[28]~q ),
	.writedata_29(\writedata[29]~q ),
	.writedata_30(\writedata[30]~q ),
	.writedata_31(\writedata[31]~q ),
	.jdo_13(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_9(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[9]~q ),
	.jdo_10(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper|the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk|jdo[10]~q ),
	.clk_clk(clk_clk));

niosLab2_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg(
	.r_sync_rst(r_sync_rst),
	.write(\write~q ),
	.address_8(\address[8]~q ),
	.address_0(\address[0]~q ),
	.address_3(\address[3]~q ),
	.address_7(\address[7]~q ),
	.address_6(\address[6]~q ),
	.address_5(\address[5]~q ),
	.address_4(\address[4]~q ),
	.address_2(\address[2]~q ),
	.address_1(\address[1]~q ),
	.debugaccess(\debugaccess~q ),
	.take_action_ocireg(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.oci_single_step_mode1(oci_single_step_mode),
	.Equal0(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.oci_ienable_16(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.oci_reg_readdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.writedata_3(\writedata[3]~q ),
	.clk_clk(clk_clk));

cyclonev_lcell_comb \read~0 (
	.dataa(!mem_used_1),
	.datab(!src_valid),
	.datac(!waitrequest),
	.datad(!src1_valid),
	.datae(!\read~q ),
	.dataf(!saved_grant_0),
	.datag(!mem),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "on";
defparam \read~0 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!mem_used_1),
	.datab(!always2),
	.datac(!waitrequest),
	.datad(!src1_valid),
	.datae(!\write~q ),
	.dataf(!saved_grant_0),
	.datag(!src_valid),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "on";
defparam \write~0 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \write~0 .shared_arith = "off";

dffeas write(
	.clk(clk_clk),
	.d(\write~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas read(
	.clk(clk_clk),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

dffeas \writedata[0] (
	.clk(clk_clk),
	.d(writedata_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[0]~q ),
	.prn(vcc));
defparam \writedata[0] .is_wysiwyg = "true";
defparam \writedata[0] .power_up = "low";

dffeas \address[3] (
	.clk(clk_clk),
	.d(address_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[3]~q ),
	.prn(vcc));
defparam \address[3] .is_wysiwyg = "true";
defparam \address[3] .power_up = "low";

dffeas \address[7] (
	.clk(clk_clk),
	.d(address_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[7]~q ),
	.prn(vcc));
defparam \address[7] .is_wysiwyg = "true";
defparam \address[7] .power_up = "low";

dffeas \address[6] (
	.clk(clk_clk),
	.d(address_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[6]~q ),
	.prn(vcc));
defparam \address[6] .is_wysiwyg = "true";
defparam \address[6] .power_up = "low";

dffeas \address[5] (
	.clk(clk_clk),
	.d(address_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[5]~q ),
	.prn(vcc));
defparam \address[5] .is_wysiwyg = "true";
defparam \address[5] .power_up = "low";

dffeas \address[4] (
	.clk(clk_clk),
	.d(address_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[4]~q ),
	.prn(vcc));
defparam \address[4] .is_wysiwyg = "true";
defparam \address[4] .power_up = "low";

dffeas \address[2] (
	.clk(clk_clk),
	.d(address_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[2]~q ),
	.prn(vcc));
defparam \address[2] .is_wysiwyg = "true";
defparam \address[2] .power_up = "low";

dffeas \address[1] (
	.clk(clk_clk),
	.d(address_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[1]~q ),
	.prn(vcc));
defparam \address[1] .is_wysiwyg = "true";
defparam \address[1] .power_up = "low";

dffeas debugaccess(
	.clk(clk_clk),
	.d(debugaccess_nxt),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\debugaccess~q ),
	.prn(vcc));
defparam debugaccess.is_wysiwyg = "true";
defparam debugaccess.power_up = "low";

dffeas \byteenable[0] (
	.clk(clk_clk),
	.d(byteenable_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[0]~q ),
	.prn(vcc));
defparam \byteenable[0] .is_wysiwyg = "true";
defparam \byteenable[0] .power_up = "low";

dffeas \writedata[1] (
	.clk(clk_clk),
	.d(writedata_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[1]~q ),
	.prn(vcc));
defparam \writedata[1] .is_wysiwyg = "true";
defparam \writedata[1] .power_up = "low";

dffeas \writedata[3] (
	.clk(clk_clk),
	.d(writedata_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[3]~q ),
	.prn(vcc));
defparam \writedata[3] .is_wysiwyg = "true";
defparam \writedata[3] .power_up = "low";

dffeas \writedata[2] (
	.clk(clk_clk),
	.d(writedata_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[2]~q ),
	.prn(vcc));
defparam \writedata[2] .is_wysiwyg = "true";
defparam \writedata[2] .power_up = "low";

dffeas \writedata[22] (
	.clk(clk_clk),
	.d(writedata_nxt[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[22]~q ),
	.prn(vcc));
defparam \writedata[22] .is_wysiwyg = "true";
defparam \writedata[22] .power_up = "low";

dffeas \byteenable[2] (
	.clk(clk_clk),
	.d(byteenable_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[2]~q ),
	.prn(vcc));
defparam \byteenable[2] .is_wysiwyg = "true";
defparam \byteenable[2] .power_up = "low";

dffeas \writedata[23] (
	.clk(clk_clk),
	.d(writedata_nxt[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[23]~q ),
	.prn(vcc));
defparam \writedata[23] .is_wysiwyg = "true";
defparam \writedata[23] .power_up = "low";

dffeas \writedata[24] (
	.clk(clk_clk),
	.d(writedata_nxt[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[24]~q ),
	.prn(vcc));
defparam \writedata[24] .is_wysiwyg = "true";
defparam \writedata[24] .power_up = "low";

dffeas \byteenable[3] (
	.clk(clk_clk),
	.d(byteenable_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[3]~q ),
	.prn(vcc));
defparam \byteenable[3] .is_wysiwyg = "true";
defparam \byteenable[3] .power_up = "low";

dffeas \writedata[25] (
	.clk(clk_clk),
	.d(writedata_nxt[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[25]~q ),
	.prn(vcc));
defparam \writedata[25] .is_wysiwyg = "true";
defparam \writedata[25] .power_up = "low";

dffeas \writedata[26] (
	.clk(clk_clk),
	.d(writedata_nxt[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[26]~q ),
	.prn(vcc));
defparam \writedata[26] .is_wysiwyg = "true";
defparam \writedata[26] .power_up = "low";

dffeas \writedata[11] (
	.clk(clk_clk),
	.d(writedata_nxt[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[11]~q ),
	.prn(vcc));
defparam \writedata[11] .is_wysiwyg = "true";
defparam \writedata[11] .power_up = "low";

dffeas \byteenable[1] (
	.clk(clk_clk),
	.d(byteenable_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[1]~q ),
	.prn(vcc));
defparam \byteenable[1] .is_wysiwyg = "true";
defparam \byteenable[1] .power_up = "low";

dffeas \writedata[12] (
	.clk(clk_clk),
	.d(writedata_nxt[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[12]~q ),
	.prn(vcc));
defparam \writedata[12] .is_wysiwyg = "true";
defparam \writedata[12] .power_up = "low";

dffeas \writedata[13] (
	.clk(clk_clk),
	.d(writedata_nxt[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[13]~q ),
	.prn(vcc));
defparam \writedata[13] .is_wysiwyg = "true";
defparam \writedata[13] .power_up = "low";

dffeas \writedata[14] (
	.clk(clk_clk),
	.d(writedata_nxt[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[14]~q ),
	.prn(vcc));
defparam \writedata[14] .is_wysiwyg = "true";
defparam \writedata[14] .power_up = "low";

dffeas \writedata[15] (
	.clk(clk_clk),
	.d(writedata_nxt[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[15]~q ),
	.prn(vcc));
defparam \writedata[15] .is_wysiwyg = "true";
defparam \writedata[15] .power_up = "low";

dffeas \writedata[16] (
	.clk(clk_clk),
	.d(writedata_nxt[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[16]~q ),
	.prn(vcc));
defparam \writedata[16] .is_wysiwyg = "true";
defparam \writedata[16] .power_up = "low";

dffeas \writedata[4] (
	.clk(clk_clk),
	.d(writedata_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[4]~q ),
	.prn(vcc));
defparam \writedata[4] .is_wysiwyg = "true";
defparam \writedata[4] .power_up = "low";

dffeas \writedata[5] (
	.clk(clk_clk),
	.d(writedata_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[5]~q ),
	.prn(vcc));
defparam \writedata[5] .is_wysiwyg = "true";
defparam \writedata[5] .power_up = "low";

dffeas \writedata[8] (
	.clk(clk_clk),
	.d(writedata_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[8]~q ),
	.prn(vcc));
defparam \writedata[8] .is_wysiwyg = "true";
defparam \writedata[8] .power_up = "low";

dffeas \writedata[10] (
	.clk(clk_clk),
	.d(writedata_nxt[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[10]~q ),
	.prn(vcc));
defparam \writedata[10] .is_wysiwyg = "true";
defparam \writedata[10] .power_up = "low";

dffeas \writedata[17] (
	.clk(clk_clk),
	.d(writedata_nxt[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[17]~q ),
	.prn(vcc));
defparam \writedata[17] .is_wysiwyg = "true";
defparam \writedata[17] .power_up = "low";

dffeas \writedata[9] (
	.clk(clk_clk),
	.d(writedata_nxt[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[9]~q ),
	.prn(vcc));
defparam \writedata[9] .is_wysiwyg = "true";
defparam \writedata[9] .power_up = "low";

dffeas \writedata[18] (
	.clk(clk_clk),
	.d(writedata_nxt[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[18]~q ),
	.prn(vcc));
defparam \writedata[18] .is_wysiwyg = "true";
defparam \writedata[18] .power_up = "low";

dffeas \writedata[19] (
	.clk(clk_clk),
	.d(writedata_nxt[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[19]~q ),
	.prn(vcc));
defparam \writedata[19] .is_wysiwyg = "true";
defparam \writedata[19] .power_up = "low";

dffeas \writedata[20] (
	.clk(clk_clk),
	.d(writedata_nxt[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[20]~q ),
	.prn(vcc));
defparam \writedata[20] .is_wysiwyg = "true";
defparam \writedata[20] .power_up = "low";

dffeas \writedata[21] (
	.clk(clk_clk),
	.d(writedata_nxt[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[21]~q ),
	.prn(vcc));
defparam \writedata[21] .is_wysiwyg = "true";
defparam \writedata[21] .power_up = "low";

dffeas \writedata[6] (
	.clk(clk_clk),
	.d(writedata_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[6]~q ),
	.prn(vcc));
defparam \writedata[6] .is_wysiwyg = "true";
defparam \writedata[6] .power_up = "low";

dffeas \writedata[7] (
	.clk(clk_clk),
	.d(writedata_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[7]~q ),
	.prn(vcc));
defparam \writedata[7] .is_wysiwyg = "true";
defparam \writedata[7] .power_up = "low";

dffeas \writedata[27] (
	.clk(clk_clk),
	.d(writedata_nxt[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[27]~q ),
	.prn(vcc));
defparam \writedata[27] .is_wysiwyg = "true";
defparam \writedata[27] .power_up = "low";

dffeas \writedata[28] (
	.clk(clk_clk),
	.d(writedata_nxt[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[28]~q ),
	.prn(vcc));
defparam \writedata[28] .is_wysiwyg = "true";
defparam \writedata[28] .power_up = "low";

dffeas \writedata[29] (
	.clk(clk_clk),
	.d(writedata_nxt[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[29]~q ),
	.prn(vcc));
defparam \writedata[29] .is_wysiwyg = "true";
defparam \writedata[29] .power_up = "low";

dffeas \writedata[30] (
	.clk(clk_clk),
	.d(writedata_nxt[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[30]~q ),
	.prn(vcc));
defparam \writedata[30] .is_wysiwyg = "true";
defparam \writedata[30] .power_up = "low";

dffeas \writedata[31] (
	.clk(clk_clk),
	.d(writedata_nxt[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[31]~q ),
	.prn(vcc));
defparam \writedata[31] .is_wysiwyg = "true";
defparam \writedata[31] .power_up = "low";

dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[22] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_22),
	.prn(vcc));
defparam \readdata[22] .is_wysiwyg = "true";
defparam \readdata[22] .power_up = "low";

dffeas \readdata[23] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_23),
	.prn(vcc));
defparam \readdata[23] .is_wysiwyg = "true";
defparam \readdata[23] .power_up = "low";

dffeas \readdata[24] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_24),
	.prn(vcc));
defparam \readdata[24] .is_wysiwyg = "true";
defparam \readdata[24] .power_up = "low";

dffeas \readdata[25] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_25),
	.prn(vcc));
defparam \readdata[25] .is_wysiwyg = "true";
defparam \readdata[25] .power_up = "low";

dffeas \readdata[26] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_26),
	.prn(vcc));
defparam \readdata[26] .is_wysiwyg = "true";
defparam \readdata[26] .power_up = "low";

dffeas \readdata[11] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

dffeas \readdata[12] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[13] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[14] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

dffeas \readdata[15] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[16] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_16),
	.prn(vcc));
defparam \readdata[16] .is_wysiwyg = "true";
defparam \readdata[16] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\readdata~1_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\readdata~2_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\readdata~3_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[17] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_17),
	.prn(vcc));
defparam \readdata[17] .is_wysiwyg = "true";
defparam \readdata[17] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[18] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_18),
	.prn(vcc));
defparam \readdata[18] .is_wysiwyg = "true";
defparam \readdata[18] .power_up = "low";

dffeas \readdata[19] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_19),
	.prn(vcc));
defparam \readdata[19] .is_wysiwyg = "true";
defparam \readdata[19] .power_up = "low";

dffeas \readdata[20] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_20),
	.prn(vcc));
defparam \readdata[20] .is_wysiwyg = "true";
defparam \readdata[20] .power_up = "low";

dffeas \readdata[21] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_21),
	.prn(vcc));
defparam \readdata[21] .is_wysiwyg = "true";
defparam \readdata[21] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[27] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_27),
	.prn(vcc));
defparam \readdata[27] .is_wysiwyg = "true";
defparam \readdata[27] .power_up = "low";

dffeas \readdata[28] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_28),
	.prn(vcc));
defparam \readdata[28] .is_wysiwyg = "true";
defparam \readdata[28] .power_up = "low";

dffeas \readdata[29] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_29),
	.prn(vcc));
defparam \readdata[29] .is_wysiwyg = "true";
defparam \readdata[29] .power_up = "low";

dffeas \readdata[30] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_30),
	.prn(vcc));
defparam \readdata[30] .is_wysiwyg = "true";
defparam \readdata[30] .power_up = "low";

dffeas \readdata[31] (
	.clk(clk_clk),
	.d(\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_31),
	.prn(vcc));
defparam \readdata[31] .is_wysiwyg = "true";
defparam \readdata[31] .power_up = "low";

dffeas \address[0] (
	.clk(clk_clk),
	.d(address_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[0]~q ),
	.prn(vcc));
defparam \address[0] .is_wysiwyg = "true";
defparam \address[0] .power_up = "low";

cyclonev_lcell_comb \readdata~0 (
	.dataa(!\address[0]~q ),
	.datab(!\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.datac(!\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug|monitor_error~q ),
	.datad(!\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~0 .extended_lut = "off";
defparam \readdata~0 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \readdata~0 .shared_arith = "off";

dffeas \address[8] (
	.clk(clk_clk),
	.d(address_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[8]~q ),
	.prn(vcc));
defparam \address[8] .is_wysiwyg = "true";
defparam \address[8] .power_up = "low";

cyclonev_lcell_comb \readdata~1 (
	.dataa(!\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug|monitor_ready~q ),
	.datab(!\address[0]~q ),
	.datac(!\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.datad(!\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~1 .extended_lut = "off";
defparam \readdata~1 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \readdata~1 .shared_arith = "off";

cyclonev_lcell_comb \readdata~2 (
	.dataa(!\address[0]~q ),
	.datab(!\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.datac(!\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datad(!\the_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug|monitor_go~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~2 .extended_lut = "off";
defparam \readdata~2 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \readdata~2 .shared_arith = "off";

cyclonev_lcell_comb \readdata~3 (
	.dataa(!\address[0]~q ),
	.datab(!\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.datac(!oci_single_step_mode),
	.datad(!\the_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~3 .extended_lut = "off";
defparam \readdata~3 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \readdata~3 .shared_arith = "off";

endmodule

module niosLab2_niosLab2_nios2_gen2_0_cpu_debug_slave_wrapper (
	break_readreg_0,
	break_readreg_1,
	MonDReg_1,
	break_readreg_2,
	MonDReg_2,
	break_readreg_3,
	MonDReg_3,
	break_readreg_16,
	MonDReg_16,
	break_readreg_24,
	MonDReg_24,
	break_readreg_4,
	break_readreg_25,
	MonDReg_25,
	break_readreg_27,
	MonDReg_27,
	break_readreg_26,
	MonDReg_26,
	MonDReg_22,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	MonDReg_23,
	MonDReg_11,
	MonDReg_13,
	MonDReg_14,
	MonDReg_10,
	MonDReg_17,
	MonDReg_9,
	MonDReg_21,
	MonDReg_6,
	break_readreg_17,
	MonDReg_7,
	break_readreg_5,
	break_readreg_28,
	MonDReg_28,
	break_readreg_29,
	MonDReg_30,
	break_readreg_30,
	break_readreg_31,
	MonDReg_31,
	break_readreg_21,
	break_readreg_18,
	break_readreg_6,
	break_readreg_22,
	break_readreg_15,
	break_readreg_23,
	break_readreg_7,
	break_readreg_13,
	break_readreg_14,
	break_readreg_10,
	break_readreg_12,
	break_readreg_11,
	break_readreg_8,
	break_readreg_9,
	sr_0,
	ir_out_0,
	ir_out_1,
	MonDReg_0,
	monitor_ready,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_1,
	ir_0,
	enable_action_strobe,
	jdo_35,
	take_action_ocimem_b,
	jdo_3,
	hbreak_enabled,
	take_action_ocimem_a,
	jdo_34,
	jdo_17,
	take_action_ocimem_a1,
	take_action_ocimem_a2,
	jdo_25,
	jdo_1,
	jdo_4,
	jdo_26,
	jdo_28,
	jdo_27,
	jdo_21,
	jdo_20,
	jdo_2,
	jdo_5,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	monitor_error,
	jdo_19,
	jdo_18,
	MonDReg_4,
	jdo_6,
	MonDReg_12,
	MonDReg_15,
	jdo_23,
	MonDReg_5,
	MonDReg_8,
	MonDReg_18,
	jdo_16,
	jdo_24,
	jdo_7,
	MonDReg_29,
	resetlatch,
	jdo_22,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_11,
	jdo_13,
	jdo_12,
	jdo_9,
	jdo_10,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	break_readreg_0;
input 	break_readreg_1;
input 	MonDReg_1;
input 	break_readreg_2;
input 	MonDReg_2;
input 	break_readreg_3;
input 	MonDReg_3;
input 	break_readreg_16;
input 	MonDReg_16;
input 	break_readreg_24;
input 	MonDReg_24;
input 	break_readreg_4;
input 	break_readreg_25;
input 	MonDReg_25;
input 	break_readreg_27;
input 	MonDReg_27;
input 	break_readreg_26;
input 	MonDReg_26;
input 	MonDReg_22;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
input 	MonDReg_23;
input 	MonDReg_11;
input 	MonDReg_13;
input 	MonDReg_14;
input 	MonDReg_10;
input 	MonDReg_17;
input 	MonDReg_9;
input 	MonDReg_21;
input 	MonDReg_6;
input 	break_readreg_17;
input 	MonDReg_7;
input 	break_readreg_5;
input 	break_readreg_28;
input 	MonDReg_28;
input 	break_readreg_29;
input 	MonDReg_30;
input 	break_readreg_30;
input 	break_readreg_31;
input 	MonDReg_31;
input 	break_readreg_21;
input 	break_readreg_18;
input 	break_readreg_6;
input 	break_readreg_22;
input 	break_readreg_15;
input 	break_readreg_23;
input 	break_readreg_7;
input 	break_readreg_13;
input 	break_readreg_14;
input 	break_readreg_10;
input 	break_readreg_12;
input 	break_readreg_11;
input 	break_readreg_8;
input 	break_readreg_9;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	MonDReg_0;
input 	monitor_ready;
output 	jdo_0;
output 	jdo_36;
output 	jdo_37;
output 	ir_1;
output 	ir_0;
output 	enable_action_strobe;
output 	jdo_35;
output 	take_action_ocimem_b;
output 	jdo_3;
input 	hbreak_enabled;
output 	take_action_ocimem_a;
output 	jdo_34;
output 	jdo_17;
output 	take_action_ocimem_a1;
output 	take_action_ocimem_a2;
output 	jdo_25;
output 	jdo_1;
output 	jdo_4;
output 	jdo_26;
output 	jdo_28;
output 	jdo_27;
output 	jdo_21;
output 	jdo_20;
output 	jdo_2;
output 	jdo_5;
output 	jdo_29;
output 	jdo_30;
output 	jdo_31;
output 	jdo_32;
output 	jdo_33;
input 	monitor_error;
output 	jdo_19;
output 	jdo_18;
input 	MonDReg_4;
output 	jdo_6;
input 	MonDReg_12;
input 	MonDReg_15;
output 	jdo_23;
input 	MonDReg_5;
input 	MonDReg_8;
input 	MonDReg_18;
output 	jdo_16;
output 	jdo_24;
output 	jdo_7;
input 	MonDReg_29;
input 	resetlatch;
output 	jdo_22;
output 	jdo_14;
output 	jdo_15;
output 	jdo_8;
output 	jdo_11;
output 	jdo_13;
output 	jdo_12;
output 	jdo_9;
output 	jdo_10;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[1]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[2]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[3]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[4]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[17]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[25]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[5]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[26]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[28]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[27]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[21]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[20]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[18]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[6]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[29]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[30]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[32]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[22]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[19]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[23]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[16]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[24]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[8]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[14]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[11]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[13]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[12]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[9]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[10]~q ;
wire \niosLab2_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_sdr~0_combout ;
wire \niosLab2_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_uir~combout ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[36]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[37]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[35]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[34]~q ;
wire \niosLab2_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_cdr~combout ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[31]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[33]~q ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[7]~q ;
wire \niosLab2_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_udr~0_combout ;
wire \the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[15]~q ;


niosLab2_niosLab2_nios2_gen2_0_cpu_debug_slave_tck the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck(
	.sr_1(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[1]~q ),
	.sr_2(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[2]~q ),
	.break_readreg_0(break_readreg_0),
	.sr_3(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[3]~q ),
	.break_readreg_1(break_readreg_1),
	.MonDReg_1(MonDReg_1),
	.sr_4(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[4]~q ),
	.break_readreg_2(break_readreg_2),
	.MonDReg_2(MonDReg_2),
	.sr_17(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[17]~q ),
	.sr_25(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[25]~q ),
	.sr_5(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[5]~q ),
	.break_readreg_3(break_readreg_3),
	.MonDReg_3(MonDReg_3),
	.sr_26(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[26]~q ),
	.sr_28(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[28]~q ),
	.sr_27(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[27]~q ),
	.sr_21(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[21]~q ),
	.sr_20(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[20]~q ),
	.sr_18(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[18]~q ),
	.break_readreg_16(break_readreg_16),
	.MonDReg_16(MonDReg_16),
	.break_readreg_24(break_readreg_24),
	.MonDReg_24(MonDReg_24),
	.sr_6(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[6]~q ),
	.break_readreg_4(break_readreg_4),
	.sr_29(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[29]~q ),
	.sr_30(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[30]~q ),
	.sr_32(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[32]~q ),
	.break_readreg_25(break_readreg_25),
	.MonDReg_25(MonDReg_25),
	.break_readreg_27(break_readreg_27),
	.MonDReg_27(MonDReg_27),
	.break_readreg_26(break_readreg_26),
	.MonDReg_26(MonDReg_26),
	.MonDReg_22(MonDReg_22),
	.sr_22(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[22]~q ),
	.break_readreg_20(break_readreg_20),
	.MonDReg_20(MonDReg_20),
	.break_readreg_19(break_readreg_19),
	.MonDReg_19(MonDReg_19),
	.sr_19(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[19]~q ),
	.MonDReg_23(MonDReg_23),
	.MonDReg_11(MonDReg_11),
	.MonDReg_13(MonDReg_13),
	.MonDReg_14(MonDReg_14),
	.MonDReg_10(MonDReg_10),
	.MonDReg_17(MonDReg_17),
	.MonDReg_9(MonDReg_9),
	.MonDReg_21(MonDReg_21),
	.MonDReg_6(MonDReg_6),
	.break_readreg_17(break_readreg_17),
	.MonDReg_7(MonDReg_7),
	.break_readreg_5(break_readreg_5),
	.break_readreg_28(break_readreg_28),
	.MonDReg_28(MonDReg_28),
	.break_readreg_29(break_readreg_29),
	.MonDReg_30(MonDReg_30),
	.break_readreg_30(break_readreg_30),
	.break_readreg_31(break_readreg_31),
	.MonDReg_31(MonDReg_31),
	.sr_23(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[23]~q ),
	.break_readreg_21(break_readreg_21),
	.break_readreg_18(break_readreg_18),
	.sr_16(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[16]~q ),
	.sr_24(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[24]~q ),
	.sr_8(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[8]~q ),
	.break_readreg_6(break_readreg_6),
	.break_readreg_22(break_readreg_22),
	.sr_14(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[14]~q ),
	.sr_11(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[11]~q ),
	.sr_13(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[13]~q ),
	.sr_12(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[12]~q ),
	.sr_9(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[9]~q ),
	.break_readreg_15(break_readreg_15),
	.sr_10(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[10]~q ),
	.break_readreg_23(break_readreg_23),
	.break_readreg_7(break_readreg_7),
	.break_readreg_13(break_readreg_13),
	.break_readreg_14(break_readreg_14),
	.break_readreg_10(break_readreg_10),
	.break_readreg_12(break_readreg_12),
	.break_readreg_11(break_readreg_11),
	.break_readreg_8(break_readreg_8),
	.break_readreg_9(break_readreg_9),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.virtual_state_sdr(\niosLab2_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_sdr~0_combout ),
	.MonDReg_0(MonDReg_0),
	.virtual_state_uir(\niosLab2_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_uir~combout ),
	.monitor_ready(monitor_ready),
	.hbreak_enabled(hbreak_enabled),
	.sr_36(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[36]~q ),
	.sr_37(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[37]~q ),
	.sr_35(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[35]~q ),
	.sr_34(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[34]~q ),
	.virtual_state_cdr(\niosLab2_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_cdr~combout ),
	.monitor_error(monitor_error),
	.MonDReg_4(MonDReg_4),
	.sr_31(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[31]~q ),
	.sr_33(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[33]~q ),
	.MonDReg_12(MonDReg_12),
	.MonDReg_15(MonDReg_15),
	.MonDReg_5(MonDReg_5),
	.MonDReg_8(MonDReg_8),
	.MonDReg_18(MonDReg_18),
	.sr_7(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[7]~q ),
	.MonDReg_29(MonDReg_29),
	.resetlatch(resetlatch),
	.sr_15(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[15]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2));

niosLab2_sld_virtual_jtag_basic_1 niosLab2_nios2_gen2_0_cpu_debug_slave_phy(
	.virtual_state_sdr(\niosLab2_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_sdr~0_combout ),
	.virtual_state_uir1(\niosLab2_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_uir~combout ),
	.virtual_state_cdr1(\niosLab2_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_cdr~combout ),
	.virtual_state_udr(\niosLab2_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_udr~0_combout ),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3));

niosLab2_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk the_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk(
	.sr_1(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[1]~q ),
	.sr_2(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[2]~q ),
	.sr_3(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[3]~q ),
	.sr_4(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[4]~q ),
	.sr_17(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[17]~q ),
	.sr_25(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[25]~q ),
	.sr_5(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[5]~q ),
	.sr_26(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[26]~q ),
	.sr_28(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[28]~q ),
	.sr_27(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[27]~q ),
	.sr_21(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[21]~q ),
	.sr_20(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[20]~q ),
	.sr_18(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[18]~q ),
	.sr_6(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[6]~q ),
	.sr_29(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[29]~q ),
	.sr_30(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[30]~q ),
	.sr_32(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[32]~q ),
	.sr_22(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[22]~q ),
	.sr_19(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[19]~q ),
	.sr_23(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[23]~q ),
	.sr_16(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[16]~q ),
	.sr_24(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[24]~q ),
	.sr_8(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[8]~q ),
	.sr_14(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[14]~q ),
	.sr_11(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[11]~q ),
	.sr_13(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[13]~q ),
	.sr_12(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[12]~q ),
	.sr_9(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[9]~q ),
	.sr_10(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[10]~q ),
	.sr_0(sr_0),
	.virtual_state_uir(\niosLab2_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_uir~combout ),
	.jdo_0(jdo_0),
	.jdo_36(jdo_36),
	.jdo_37(jdo_37),
	.ir_1(ir_1),
	.ir_0(ir_0),
	.enable_action_strobe1(enable_action_strobe),
	.jdo_35(jdo_35),
	.take_action_ocimem_b1(take_action_ocimem_b),
	.jdo_3(jdo_3),
	.take_action_ocimem_a1(take_action_ocimem_a),
	.jdo_34(jdo_34),
	.jdo_17(jdo_17),
	.take_action_ocimem_a2(take_action_ocimem_a1),
	.take_action_ocimem_a3(take_action_ocimem_a2),
	.jdo_25(jdo_25),
	.jdo_1(jdo_1),
	.jdo_4(jdo_4),
	.sr_36(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[36]~q ),
	.sr_37(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[37]~q ),
	.sr_35(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[35]~q ),
	.jdo_26(jdo_26),
	.jdo_28(jdo_28),
	.jdo_27(jdo_27),
	.jdo_21(jdo_21),
	.jdo_20(jdo_20),
	.sr_34(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[34]~q ),
	.jdo_2(jdo_2),
	.jdo_5(jdo_5),
	.jdo_29(jdo_29),
	.jdo_30(jdo_30),
	.jdo_31(jdo_31),
	.jdo_32(jdo_32),
	.jdo_33(jdo_33),
	.jdo_19(jdo_19),
	.jdo_18(jdo_18),
	.jdo_6(jdo_6),
	.sr_31(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[31]~q ),
	.sr_33(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[33]~q ),
	.jdo_23(jdo_23),
	.jdo_16(jdo_16),
	.jdo_24(jdo_24),
	.sr_7(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[7]~q ),
	.jdo_7(jdo_7),
	.virtual_state_udr(\niosLab2_nios2_gen2_0_cpu_debug_slave_phy|virtual_state_udr~0_combout ),
	.jdo_22(jdo_22),
	.jdo_14(jdo_14),
	.jdo_15(jdo_15),
	.jdo_8(jdo_8),
	.jdo_11(jdo_11),
	.jdo_13(jdo_13),
	.jdo_12(jdo_12),
	.jdo_9(jdo_9),
	.jdo_10(jdo_10),
	.sr_15(\the_niosLab2_nios2_gen2_0_cpu_debug_slave_tck|sr[15]~q ),
	.ir_in({irf_reg_1_2,irf_reg_0_2}),
	.clk_clk(clk_clk));

endmodule

module niosLab2_niosLab2_nios2_gen2_0_cpu_debug_slave_sysclk (
	sr_1,
	sr_2,
	sr_3,
	sr_4,
	sr_17,
	sr_25,
	sr_5,
	sr_26,
	sr_28,
	sr_27,
	sr_21,
	sr_20,
	sr_18,
	sr_6,
	sr_29,
	sr_30,
	sr_32,
	sr_22,
	sr_19,
	sr_23,
	sr_16,
	sr_24,
	sr_8,
	sr_14,
	sr_11,
	sr_13,
	sr_12,
	sr_9,
	sr_10,
	sr_0,
	virtual_state_uir,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_1,
	ir_0,
	enable_action_strobe1,
	jdo_35,
	take_action_ocimem_b1,
	jdo_3,
	take_action_ocimem_a1,
	jdo_34,
	jdo_17,
	take_action_ocimem_a2,
	take_action_ocimem_a3,
	jdo_25,
	jdo_1,
	jdo_4,
	sr_36,
	sr_37,
	sr_35,
	jdo_26,
	jdo_28,
	jdo_27,
	jdo_21,
	jdo_20,
	sr_34,
	jdo_2,
	jdo_5,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	jdo_19,
	jdo_18,
	jdo_6,
	sr_31,
	sr_33,
	jdo_23,
	jdo_16,
	jdo_24,
	sr_7,
	jdo_7,
	virtual_state_udr,
	jdo_22,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_11,
	jdo_13,
	jdo_12,
	jdo_9,
	jdo_10,
	sr_15,
	ir_in,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	sr_1;
input 	sr_2;
input 	sr_3;
input 	sr_4;
input 	sr_17;
input 	sr_25;
input 	sr_5;
input 	sr_26;
input 	sr_28;
input 	sr_27;
input 	sr_21;
input 	sr_20;
input 	sr_18;
input 	sr_6;
input 	sr_29;
input 	sr_30;
input 	sr_32;
input 	sr_22;
input 	sr_19;
input 	sr_23;
input 	sr_16;
input 	sr_24;
input 	sr_8;
input 	sr_14;
input 	sr_11;
input 	sr_13;
input 	sr_12;
input 	sr_9;
input 	sr_10;
input 	sr_0;
input 	virtual_state_uir;
output 	jdo_0;
output 	jdo_36;
output 	jdo_37;
output 	ir_1;
output 	ir_0;
output 	enable_action_strobe1;
output 	jdo_35;
output 	take_action_ocimem_b1;
output 	jdo_3;
output 	take_action_ocimem_a1;
output 	jdo_34;
output 	jdo_17;
output 	take_action_ocimem_a2;
output 	take_action_ocimem_a3;
output 	jdo_25;
output 	jdo_1;
output 	jdo_4;
input 	sr_36;
input 	sr_37;
input 	sr_35;
output 	jdo_26;
output 	jdo_28;
output 	jdo_27;
output 	jdo_21;
output 	jdo_20;
input 	sr_34;
output 	jdo_2;
output 	jdo_5;
output 	jdo_29;
output 	jdo_30;
output 	jdo_31;
output 	jdo_32;
output 	jdo_33;
output 	jdo_19;
output 	jdo_18;
output 	jdo_6;
input 	sr_31;
input 	sr_33;
output 	jdo_23;
output 	jdo_16;
output 	jdo_24;
input 	sr_7;
output 	jdo_7;
input 	virtual_state_udr;
output 	jdo_22;
output 	jdo_14;
output 	jdo_15;
output 	jdo_8;
output 	jdo_11;
output 	jdo_13;
output 	jdo_12;
output 	jdo_9;
output 	jdo_10;
input 	sr_15;
input 	[1:0] ir_in;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer3|dreg[0]~q ;
wire \the_altera_std_synchronizer4|dreg[0]~q ;
wire \sync2_udr~q ;
wire \update_jdo_strobe~0_combout ;
wire \update_jdo_strobe~q ;
wire \sync2_uir~q ;
wire \jxuir~0_combout ;
wire \jxuir~q ;


niosLab2_altera_std_synchronizer_1 the_altera_std_synchronizer4(
	.din(virtual_state_uir),
	.dreg_0(\the_altera_std_synchronizer4|dreg[0]~q ),
	.clk(clk_clk));

niosLab2_altera_std_synchronizer the_altera_std_synchronizer3(
	.dreg_0(\the_altera_std_synchronizer3|dreg[0]~q ),
	.din(virtual_state_udr),
	.clk(clk_clk));

dffeas \jdo[0] (
	.clk(clk_clk),
	.d(sr_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_0),
	.prn(vcc));
defparam \jdo[0] .is_wysiwyg = "true";
defparam \jdo[0] .power_up = "low";

dffeas \jdo[36] (
	.clk(clk_clk),
	.d(sr_36),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_36),
	.prn(vcc));
defparam \jdo[36] .is_wysiwyg = "true";
defparam \jdo[36] .power_up = "low";

dffeas \jdo[37] (
	.clk(clk_clk),
	.d(sr_37),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_37),
	.prn(vcc));
defparam \jdo[37] .is_wysiwyg = "true";
defparam \jdo[37] .power_up = "low";

dffeas \ir[1] (
	.clk(clk_clk),
	.d(ir_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(ir_1),
	.prn(vcc));
defparam \ir[1] .is_wysiwyg = "true";
defparam \ir[1] .power_up = "low";

dffeas \ir[0] (
	.clk(clk_clk),
	.d(ir_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(ir_0),
	.prn(vcc));
defparam \ir[0] .is_wysiwyg = "true";
defparam \ir[0] .power_up = "low";

dffeas enable_action_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(enable_action_strobe1),
	.prn(vcc));
defparam enable_action_strobe.is_wysiwyg = "true";
defparam enable_action_strobe.power_up = "low";

dffeas \jdo[35] (
	.clk(clk_clk),
	.d(sr_35),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_35),
	.prn(vcc));
defparam \jdo[35] .is_wysiwyg = "true";
defparam \jdo[35] .power_up = "low";

cyclonev_lcell_comb take_action_ocimem_b(
	.dataa(!ir_1),
	.datab(!ir_0),
	.datac(!enable_action_strobe1),
	.datad(!jdo_35),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_b1),
	.sumout(),
	.cout(),
	.shareout());
defparam take_action_ocimem_b.extended_lut = "off";
defparam take_action_ocimem_b.lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam take_action_ocimem_b.shared_arith = "off";

dffeas \jdo[3] (
	.clk(clk_clk),
	.d(sr_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_3),
	.prn(vcc));
defparam \jdo[3] .is_wysiwyg = "true";
defparam \jdo[3] .power_up = "low";

cyclonev_lcell_comb \take_action_ocimem_a~0 (
	.dataa(!ir_1),
	.datab(!ir_0),
	.datac(!enable_action_strobe1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_a1),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_ocimem_a~0 .extended_lut = "off";
defparam \take_action_ocimem_a~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \take_action_ocimem_a~0 .shared_arith = "off";

dffeas \jdo[34] (
	.clk(clk_clk),
	.d(sr_34),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_34),
	.prn(vcc));
defparam \jdo[34] .is_wysiwyg = "true";
defparam \jdo[34] .power_up = "low";

dffeas \jdo[17] (
	.clk(clk_clk),
	.d(sr_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_17),
	.prn(vcc));
defparam \jdo[17] .is_wysiwyg = "true";
defparam \jdo[17] .power_up = "low";

cyclonev_lcell_comb \take_action_ocimem_a~1 (
	.dataa(!ir_1),
	.datab(!ir_0),
	.datac(!enable_action_strobe1),
	.datad(!jdo_35),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_a2),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_ocimem_a~1 .extended_lut = "off";
defparam \take_action_ocimem_a~1 .lut_mask = 64'hFFEFFFEFFFEFFFEF;
defparam \take_action_ocimem_a~1 .shared_arith = "off";

cyclonev_lcell_comb take_action_ocimem_a(
	.dataa(!take_action_ocimem_a2),
	.datab(!jdo_34),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_a3),
	.sumout(),
	.cout(),
	.shareout());
defparam take_action_ocimem_a.extended_lut = "off";
defparam take_action_ocimem_a.lut_mask = 64'h7777777777777777;
defparam take_action_ocimem_a.shared_arith = "off";

dffeas \jdo[25] (
	.clk(clk_clk),
	.d(sr_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_25),
	.prn(vcc));
defparam \jdo[25] .is_wysiwyg = "true";
defparam \jdo[25] .power_up = "low";

dffeas \jdo[1] (
	.clk(clk_clk),
	.d(sr_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_1),
	.prn(vcc));
defparam \jdo[1] .is_wysiwyg = "true";
defparam \jdo[1] .power_up = "low";

dffeas \jdo[4] (
	.clk(clk_clk),
	.d(sr_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_4),
	.prn(vcc));
defparam \jdo[4] .is_wysiwyg = "true";
defparam \jdo[4] .power_up = "low";

dffeas \jdo[26] (
	.clk(clk_clk),
	.d(sr_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_26),
	.prn(vcc));
defparam \jdo[26] .is_wysiwyg = "true";
defparam \jdo[26] .power_up = "low";

dffeas \jdo[28] (
	.clk(clk_clk),
	.d(sr_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_28),
	.prn(vcc));
defparam \jdo[28] .is_wysiwyg = "true";
defparam \jdo[28] .power_up = "low";

dffeas \jdo[27] (
	.clk(clk_clk),
	.d(sr_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_27),
	.prn(vcc));
defparam \jdo[27] .is_wysiwyg = "true";
defparam \jdo[27] .power_up = "low";

dffeas \jdo[21] (
	.clk(clk_clk),
	.d(sr_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_21),
	.prn(vcc));
defparam \jdo[21] .is_wysiwyg = "true";
defparam \jdo[21] .power_up = "low";

dffeas \jdo[20] (
	.clk(clk_clk),
	.d(sr_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_20),
	.prn(vcc));
defparam \jdo[20] .is_wysiwyg = "true";
defparam \jdo[20] .power_up = "low";

dffeas \jdo[2] (
	.clk(clk_clk),
	.d(sr_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_2),
	.prn(vcc));
defparam \jdo[2] .is_wysiwyg = "true";
defparam \jdo[2] .power_up = "low";

dffeas \jdo[5] (
	.clk(clk_clk),
	.d(sr_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_5),
	.prn(vcc));
defparam \jdo[5] .is_wysiwyg = "true";
defparam \jdo[5] .power_up = "low";

dffeas \jdo[29] (
	.clk(clk_clk),
	.d(sr_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_29),
	.prn(vcc));
defparam \jdo[29] .is_wysiwyg = "true";
defparam \jdo[29] .power_up = "low";

dffeas \jdo[30] (
	.clk(clk_clk),
	.d(sr_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_30),
	.prn(vcc));
defparam \jdo[30] .is_wysiwyg = "true";
defparam \jdo[30] .power_up = "low";

dffeas \jdo[31] (
	.clk(clk_clk),
	.d(sr_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_31),
	.prn(vcc));
defparam \jdo[31] .is_wysiwyg = "true";
defparam \jdo[31] .power_up = "low";

dffeas \jdo[32] (
	.clk(clk_clk),
	.d(sr_32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_32),
	.prn(vcc));
defparam \jdo[32] .is_wysiwyg = "true";
defparam \jdo[32] .power_up = "low";

dffeas \jdo[33] (
	.clk(clk_clk),
	.d(sr_33),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_33),
	.prn(vcc));
defparam \jdo[33] .is_wysiwyg = "true";
defparam \jdo[33] .power_up = "low";

dffeas \jdo[19] (
	.clk(clk_clk),
	.d(sr_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_19),
	.prn(vcc));
defparam \jdo[19] .is_wysiwyg = "true";
defparam \jdo[19] .power_up = "low";

dffeas \jdo[18] (
	.clk(clk_clk),
	.d(sr_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_18),
	.prn(vcc));
defparam \jdo[18] .is_wysiwyg = "true";
defparam \jdo[18] .power_up = "low";

dffeas \jdo[6] (
	.clk(clk_clk),
	.d(sr_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_6),
	.prn(vcc));
defparam \jdo[6] .is_wysiwyg = "true";
defparam \jdo[6] .power_up = "low";

dffeas \jdo[23] (
	.clk(clk_clk),
	.d(sr_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_23),
	.prn(vcc));
defparam \jdo[23] .is_wysiwyg = "true";
defparam \jdo[23] .power_up = "low";

dffeas \jdo[16] (
	.clk(clk_clk),
	.d(sr_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_16),
	.prn(vcc));
defparam \jdo[16] .is_wysiwyg = "true";
defparam \jdo[16] .power_up = "low";

dffeas \jdo[24] (
	.clk(clk_clk),
	.d(sr_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_24),
	.prn(vcc));
defparam \jdo[24] .is_wysiwyg = "true";
defparam \jdo[24] .power_up = "low";

dffeas \jdo[7] (
	.clk(clk_clk),
	.d(sr_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_7),
	.prn(vcc));
defparam \jdo[7] .is_wysiwyg = "true";
defparam \jdo[7] .power_up = "low";

dffeas \jdo[22] (
	.clk(clk_clk),
	.d(sr_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_22),
	.prn(vcc));
defparam \jdo[22] .is_wysiwyg = "true";
defparam \jdo[22] .power_up = "low";

dffeas \jdo[14] (
	.clk(clk_clk),
	.d(sr_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_14),
	.prn(vcc));
defparam \jdo[14] .is_wysiwyg = "true";
defparam \jdo[14] .power_up = "low";

dffeas \jdo[15] (
	.clk(clk_clk),
	.d(sr_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_15),
	.prn(vcc));
defparam \jdo[15] .is_wysiwyg = "true";
defparam \jdo[15] .power_up = "low";

dffeas \jdo[8] (
	.clk(clk_clk),
	.d(sr_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_8),
	.prn(vcc));
defparam \jdo[8] .is_wysiwyg = "true";
defparam \jdo[8] .power_up = "low";

dffeas \jdo[11] (
	.clk(clk_clk),
	.d(sr_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_11),
	.prn(vcc));
defparam \jdo[11] .is_wysiwyg = "true";
defparam \jdo[11] .power_up = "low";

dffeas \jdo[13] (
	.clk(clk_clk),
	.d(sr_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_13),
	.prn(vcc));
defparam \jdo[13] .is_wysiwyg = "true";
defparam \jdo[13] .power_up = "low";

dffeas \jdo[12] (
	.clk(clk_clk),
	.d(sr_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_12),
	.prn(vcc));
defparam \jdo[12] .is_wysiwyg = "true";
defparam \jdo[12] .power_up = "low";

dffeas \jdo[9] (
	.clk(clk_clk),
	.d(sr_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_9),
	.prn(vcc));
defparam \jdo[9] .is_wysiwyg = "true";
defparam \jdo[9] .power_up = "low";

dffeas \jdo[10] (
	.clk(clk_clk),
	.d(sr_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_10),
	.prn(vcc));
defparam \jdo[10] .is_wysiwyg = "true";
defparam \jdo[10] .power_up = "low";

dffeas sync2_udr(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer3|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_udr~q ),
	.prn(vcc));
defparam sync2_udr.is_wysiwyg = "true";
defparam sync2_udr.power_up = "low";

cyclonev_lcell_comb \update_jdo_strobe~0 (
	.dataa(!\sync2_udr~q ),
	.datab(!\the_altera_std_synchronizer3|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_jdo_strobe~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_jdo_strobe~0 .extended_lut = "off";
defparam \update_jdo_strobe~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \update_jdo_strobe~0 .shared_arith = "off";

dffeas update_jdo_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\update_jdo_strobe~q ),
	.prn(vcc));
defparam update_jdo_strobe.is_wysiwyg = "true";
defparam update_jdo_strobe.power_up = "low";

dffeas sync2_uir(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer4|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_uir~q ),
	.prn(vcc));
defparam sync2_uir.is_wysiwyg = "true";
defparam sync2_uir.power_up = "low";

cyclonev_lcell_comb \jxuir~0 (
	.dataa(!\sync2_uir~q ),
	.datab(!\the_altera_std_synchronizer4|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jxuir~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jxuir~0 .extended_lut = "off";
defparam \jxuir~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \jxuir~0 .shared_arith = "off";

dffeas jxuir(
	.clk(clk_clk),
	.d(\jxuir~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jxuir~q ),
	.prn(vcc));
defparam jxuir.is_wysiwyg = "true";
defparam jxuir.power_up = "low";

endmodule

module niosLab2_altera_std_synchronizer (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosLab2_altera_std_synchronizer_1 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosLab2_niosLab2_nios2_gen2_0_cpu_debug_slave_tck (
	sr_1,
	sr_2,
	break_readreg_0,
	sr_3,
	break_readreg_1,
	MonDReg_1,
	sr_4,
	break_readreg_2,
	MonDReg_2,
	sr_17,
	sr_25,
	sr_5,
	break_readreg_3,
	MonDReg_3,
	sr_26,
	sr_28,
	sr_27,
	sr_21,
	sr_20,
	sr_18,
	break_readreg_16,
	MonDReg_16,
	break_readreg_24,
	MonDReg_24,
	sr_6,
	break_readreg_4,
	sr_29,
	sr_30,
	sr_32,
	break_readreg_25,
	MonDReg_25,
	break_readreg_27,
	MonDReg_27,
	break_readreg_26,
	MonDReg_26,
	MonDReg_22,
	sr_22,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	sr_19,
	MonDReg_23,
	MonDReg_11,
	MonDReg_13,
	MonDReg_14,
	MonDReg_10,
	MonDReg_17,
	MonDReg_9,
	MonDReg_21,
	MonDReg_6,
	break_readreg_17,
	MonDReg_7,
	break_readreg_5,
	break_readreg_28,
	MonDReg_28,
	break_readreg_29,
	MonDReg_30,
	break_readreg_30,
	break_readreg_31,
	MonDReg_31,
	sr_23,
	break_readreg_21,
	break_readreg_18,
	sr_16,
	sr_24,
	sr_8,
	break_readreg_6,
	break_readreg_22,
	sr_14,
	sr_11,
	sr_13,
	sr_12,
	sr_9,
	break_readreg_15,
	sr_10,
	break_readreg_23,
	break_readreg_7,
	break_readreg_13,
	break_readreg_14,
	break_readreg_10,
	break_readreg_12,
	break_readreg_11,
	break_readreg_8,
	break_readreg_9,
	sr_0,
	ir_out_0,
	ir_out_1,
	virtual_state_sdr,
	MonDReg_0,
	virtual_state_uir,
	monitor_ready,
	hbreak_enabled,
	sr_36,
	sr_37,
	sr_35,
	sr_34,
	virtual_state_cdr,
	monitor_error,
	MonDReg_4,
	sr_31,
	sr_33,
	MonDReg_12,
	MonDReg_15,
	MonDReg_5,
	MonDReg_8,
	MonDReg_18,
	sr_7,
	MonDReg_29,
	resetlatch,
	sr_15,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2)/* synthesis synthesis_greybox=1 */;
output 	sr_1;
output 	sr_2;
input 	break_readreg_0;
output 	sr_3;
input 	break_readreg_1;
input 	MonDReg_1;
output 	sr_4;
input 	break_readreg_2;
input 	MonDReg_2;
output 	sr_17;
output 	sr_25;
output 	sr_5;
input 	break_readreg_3;
input 	MonDReg_3;
output 	sr_26;
output 	sr_28;
output 	sr_27;
output 	sr_21;
output 	sr_20;
output 	sr_18;
input 	break_readreg_16;
input 	MonDReg_16;
input 	break_readreg_24;
input 	MonDReg_24;
output 	sr_6;
input 	break_readreg_4;
output 	sr_29;
output 	sr_30;
output 	sr_32;
input 	break_readreg_25;
input 	MonDReg_25;
input 	break_readreg_27;
input 	MonDReg_27;
input 	break_readreg_26;
input 	MonDReg_26;
input 	MonDReg_22;
output 	sr_22;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
output 	sr_19;
input 	MonDReg_23;
input 	MonDReg_11;
input 	MonDReg_13;
input 	MonDReg_14;
input 	MonDReg_10;
input 	MonDReg_17;
input 	MonDReg_9;
input 	MonDReg_21;
input 	MonDReg_6;
input 	break_readreg_17;
input 	MonDReg_7;
input 	break_readreg_5;
input 	break_readreg_28;
input 	MonDReg_28;
input 	break_readreg_29;
input 	MonDReg_30;
input 	break_readreg_30;
input 	break_readreg_31;
input 	MonDReg_31;
output 	sr_23;
input 	break_readreg_21;
input 	break_readreg_18;
output 	sr_16;
output 	sr_24;
output 	sr_8;
input 	break_readreg_6;
input 	break_readreg_22;
output 	sr_14;
output 	sr_11;
output 	sr_13;
output 	sr_12;
output 	sr_9;
input 	break_readreg_15;
output 	sr_10;
input 	break_readreg_23;
input 	break_readreg_7;
input 	break_readreg_13;
input 	break_readreg_14;
input 	break_readreg_10;
input 	break_readreg_12;
input 	break_readreg_11;
input 	break_readreg_8;
input 	break_readreg_9;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	virtual_state_sdr;
input 	MonDReg_0;
input 	virtual_state_uir;
input 	monitor_ready;
input 	hbreak_enabled;
output 	sr_36;
output 	sr_37;
output 	sr_35;
output 	sr_34;
input 	virtual_state_cdr;
input 	monitor_error;
input 	MonDReg_4;
output 	sr_31;
output 	sr_33;
input 	MonDReg_12;
input 	MonDReg_15;
input 	MonDReg_5;
input 	MonDReg_8;
input 	MonDReg_18;
output 	sr_7;
input 	MonDReg_29;
input 	resetlatch;
output 	sr_15;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer2|dreg[0]~q ;
wire \the_altera_std_synchronizer1|dreg[0]~q ;
wire \sr~8_combout ;
wire \sr[14]~9_combout ;
wire \sr[14]~10_combout ;
wire \sr~11_combout ;
wire \sr~12_combout ;
wire \sr~13_combout ;
wire \sr~20_combout ;
wire \sr[29]~21_combout ;
wire \sr[29]~19_combout ;
wire \sr~22_combout ;
wire \sr~23_combout ;
wire \sr~24_combout ;
wire \sr~25_combout ;
wire \sr~26_combout ;
wire \sr~27_combout ;
wire \sr~28_combout ;
wire \sr~29_combout ;
wire \sr~30_combout ;
wire \sr~31_combout ;
wire \sr~32_combout ;
wire \sr~37_combout ;
wire \sr~39_combout ;
wire \sr~40_combout ;
wire \sr~43_combout ;
wire \sr~44_combout ;
wire \sr~45_combout ;
wire \sr~46_combout ;
wire \sr~47_combout ;
wire \sr~50_combout ;
wire \sr~51_combout ;
wire \sr~52_combout ;
wire \sr~53_combout ;
wire \sr~54_combout ;
wire \sr~5_combout ;
wire \sr~6_combout ;
wire \DRsize.000~q ;
wire \sr~7_combout ;
wire \sr~14_combout ;
wire \sr[37]~15_combout ;
wire \sr~16_combout ;
wire \Mux37~0_combout ;
wire \DRsize.100~q ;
wire \sr~56_combout ;
wire \sr~17_combout ;
wire \sr~18_combout ;
wire \sr[29]~33_combout ;
wire \sr~34_combout ;
wire \sr~35_combout ;
wire \sr~36_combout ;
wire \sr~38_combout ;
wire \sr~41_combout ;
wire \sr~42_combout ;
wire \sr[29]~55_combout ;
wire \DRsize.010~q ;
wire \sr~48_combout ;
wire \sr~49_combout ;


niosLab2_altera_std_synchronizer_3 the_altera_std_synchronizer2(
	.dreg_0(\the_altera_std_synchronizer2|dreg[0]~q ),
	.din(monitor_ready),
	.clk(altera_internal_jtag));

niosLab2_altera_std_synchronizer_2 the_altera_std_synchronizer1(
	.dreg_0(\the_altera_std_synchronizer1|dreg[0]~q ),
	.din(hbreak_enabled),
	.clk(altera_internal_jtag));

dffeas \sr[1] (
	.clk(altera_internal_jtag),
	.d(\sr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_1),
	.prn(vcc));
defparam \sr[1] .is_wysiwyg = "true";
defparam \sr[1] .power_up = "low";

dffeas \sr[2] (
	.clk(altera_internal_jtag),
	.d(\sr~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_2),
	.prn(vcc));
defparam \sr[2] .is_wysiwyg = "true";
defparam \sr[2] .power_up = "low";

dffeas \sr[3] (
	.clk(altera_internal_jtag),
	.d(\sr~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_3),
	.prn(vcc));
defparam \sr[3] .is_wysiwyg = "true";
defparam \sr[3] .power_up = "low";

dffeas \sr[4] (
	.clk(altera_internal_jtag),
	.d(\sr~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_4),
	.prn(vcc));
defparam \sr[4] .is_wysiwyg = "true";
defparam \sr[4] .power_up = "low";

dffeas \sr[17] (
	.clk(altera_internal_jtag),
	.d(\sr~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~21_combout ),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_17),
	.prn(vcc));
defparam \sr[17] .is_wysiwyg = "true";
defparam \sr[17] .power_up = "low";

dffeas \sr[25] (
	.clk(altera_internal_jtag),
	.d(\sr~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~21_combout ),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_25),
	.prn(vcc));
defparam \sr[25] .is_wysiwyg = "true";
defparam \sr[25] .power_up = "low";

dffeas \sr[5] (
	.clk(altera_internal_jtag),
	.d(\sr~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_5),
	.prn(vcc));
defparam \sr[5] .is_wysiwyg = "true";
defparam \sr[5] .power_up = "low";

dffeas \sr[26] (
	.clk(altera_internal_jtag),
	.d(\sr~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~21_combout ),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_26),
	.prn(vcc));
defparam \sr[26] .is_wysiwyg = "true";
defparam \sr[26] .power_up = "low";

dffeas \sr[28] (
	.clk(altera_internal_jtag),
	.d(\sr~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~21_combout ),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_28),
	.prn(vcc));
defparam \sr[28] .is_wysiwyg = "true";
defparam \sr[28] .power_up = "low";

dffeas \sr[27] (
	.clk(altera_internal_jtag),
	.d(\sr~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~21_combout ),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_27),
	.prn(vcc));
defparam \sr[27] .is_wysiwyg = "true";
defparam \sr[27] .power_up = "low";

dffeas \sr[21] (
	.clk(altera_internal_jtag),
	.d(\sr~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~21_combout ),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_21),
	.prn(vcc));
defparam \sr[21] .is_wysiwyg = "true";
defparam \sr[21] .power_up = "low";

dffeas \sr[20] (
	.clk(altera_internal_jtag),
	.d(\sr~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~21_combout ),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_20),
	.prn(vcc));
defparam \sr[20] .is_wysiwyg = "true";
defparam \sr[20] .power_up = "low";

dffeas \sr[18] (
	.clk(altera_internal_jtag),
	.d(\sr~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~21_combout ),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_18),
	.prn(vcc));
defparam \sr[18] .is_wysiwyg = "true";
defparam \sr[18] .power_up = "low";

dffeas \sr[6] (
	.clk(altera_internal_jtag),
	.d(\sr~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_6),
	.prn(vcc));
defparam \sr[6] .is_wysiwyg = "true";
defparam \sr[6] .power_up = "low";

dffeas \sr[29] (
	.clk(altera_internal_jtag),
	.d(\sr~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~21_combout ),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_29),
	.prn(vcc));
defparam \sr[29] .is_wysiwyg = "true";
defparam \sr[29] .power_up = "low";

dffeas \sr[30] (
	.clk(altera_internal_jtag),
	.d(\sr~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~21_combout ),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_30),
	.prn(vcc));
defparam \sr[30] .is_wysiwyg = "true";
defparam \sr[30] .power_up = "low";

dffeas \sr[32] (
	.clk(altera_internal_jtag),
	.d(\sr~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~21_combout ),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_32),
	.prn(vcc));
defparam \sr[32] .is_wysiwyg = "true";
defparam \sr[32] .power_up = "low";

dffeas \sr[22] (
	.clk(altera_internal_jtag),
	.d(\sr~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~21_combout ),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_22),
	.prn(vcc));
defparam \sr[22] .is_wysiwyg = "true";
defparam \sr[22] .power_up = "low";

dffeas \sr[19] (
	.clk(altera_internal_jtag),
	.d(\sr~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~21_combout ),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_19),
	.prn(vcc));
defparam \sr[19] .is_wysiwyg = "true";
defparam \sr[19] .power_up = "low";

dffeas \sr[23] (
	.clk(altera_internal_jtag),
	.d(\sr~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~21_combout ),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_23),
	.prn(vcc));
defparam \sr[23] .is_wysiwyg = "true";
defparam \sr[23] .power_up = "low";

dffeas \sr[16] (
	.clk(altera_internal_jtag),
	.d(\sr~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~21_combout ),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_16),
	.prn(vcc));
defparam \sr[16] .is_wysiwyg = "true";
defparam \sr[16] .power_up = "low";

dffeas \sr[24] (
	.clk(altera_internal_jtag),
	.d(\sr~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~21_combout ),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_24),
	.prn(vcc));
defparam \sr[24] .is_wysiwyg = "true";
defparam \sr[24] .power_up = "low";

dffeas \sr[8] (
	.clk(altera_internal_jtag),
	.d(\sr~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_8),
	.prn(vcc));
defparam \sr[8] .is_wysiwyg = "true";
defparam \sr[8] .power_up = "low";

dffeas \sr[14] (
	.clk(altera_internal_jtag),
	.d(\sr~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_14),
	.prn(vcc));
defparam \sr[14] .is_wysiwyg = "true";
defparam \sr[14] .power_up = "low";

dffeas \sr[11] (
	.clk(altera_internal_jtag),
	.d(\sr~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_11),
	.prn(vcc));
defparam \sr[11] .is_wysiwyg = "true";
defparam \sr[11] .power_up = "low";

dffeas \sr[13] (
	.clk(altera_internal_jtag),
	.d(\sr~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_13),
	.prn(vcc));
defparam \sr[13] .is_wysiwyg = "true";
defparam \sr[13] .power_up = "low";

dffeas \sr[12] (
	.clk(altera_internal_jtag),
	.d(\sr~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_12),
	.prn(vcc));
defparam \sr[12] .is_wysiwyg = "true";
defparam \sr[12] .power_up = "low";

dffeas \sr[9] (
	.clk(altera_internal_jtag),
	.d(\sr~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_9),
	.prn(vcc));
defparam \sr[9] .is_wysiwyg = "true";
defparam \sr[9] .power_up = "low";

dffeas \sr[10] (
	.clk(altera_internal_jtag),
	.d(\sr~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[14]~9_combout ),
	.sload(gnd),
	.ena(\sr[14]~10_combout ),
	.q(sr_10),
	.prn(vcc));
defparam \sr[10] .is_wysiwyg = "true";
defparam \sr[10] .power_up = "low";

dffeas \sr[0] (
	.clk(altera_internal_jtag),
	.d(\sr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_0),
	.prn(vcc));
defparam \sr[0] .is_wysiwyg = "true";
defparam \sr[0] .power_up = "low";

dffeas \ir_out[0] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer2|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_0),
	.prn(vcc));
defparam \ir_out[0] .is_wysiwyg = "true";
defparam \ir_out[0] .power_up = "low";

dffeas \ir_out[1] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer1|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_1),
	.prn(vcc));
defparam \ir_out[1] .is_wysiwyg = "true";
defparam \ir_out[1] .power_up = "low";

dffeas \sr[36] (
	.clk(altera_internal_jtag),
	.d(\sr~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[37]~15_combout ),
	.q(sr_36),
	.prn(vcc));
defparam \sr[36] .is_wysiwyg = "true";
defparam \sr[36] .power_up = "low";

dffeas \sr[37] (
	.clk(altera_internal_jtag),
	.d(\sr~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[37]~15_combout ),
	.q(sr_37),
	.prn(vcc));
defparam \sr[37] .is_wysiwyg = "true";
defparam \sr[37] .power_up = "low";

dffeas \sr[35] (
	.clk(altera_internal_jtag),
	.d(\sr~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_35),
	.prn(vcc));
defparam \sr[35] .is_wysiwyg = "true";
defparam \sr[35] .power_up = "low";

dffeas \sr[34] (
	.clk(altera_internal_jtag),
	.d(\sr~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_34),
	.prn(vcc));
defparam \sr[34] .is_wysiwyg = "true";
defparam \sr[34] .power_up = "low";

dffeas \sr[31] (
	.clk(altera_internal_jtag),
	.d(\sr~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_31),
	.prn(vcc));
defparam \sr[31] .is_wysiwyg = "true";
defparam \sr[31] .power_up = "low";

dffeas \sr[33] (
	.clk(altera_internal_jtag),
	.d(\sr~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~19_combout ),
	.q(sr_33),
	.prn(vcc));
defparam \sr[33] .is_wysiwyg = "true";
defparam \sr[33] .power_up = "low";

dffeas \sr[7] (
	.clk(altera_internal_jtag),
	.d(\sr~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_7),
	.prn(vcc));
defparam \sr[7] .is_wysiwyg = "true";
defparam \sr[7] .power_up = "low";

dffeas \sr[15] (
	.clk(altera_internal_jtag),
	.d(\sr~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_15),
	.prn(vcc));
defparam \sr[15] .is_wysiwyg = "true";
defparam \sr[15] .power_up = "low";

cyclonev_lcell_comb \sr~8 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_2),
	.datad(!break_readreg_0),
	.datae(!MonDReg_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~8 .extended_lut = "off";
defparam \sr~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~8 .shared_arith = "off";

cyclonev_lcell_comb \sr[14]~9 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!irf_reg_0_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[14]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[14]~9 .extended_lut = "off";
defparam \sr[14]~9 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \sr[14]~9 .shared_arith = "off";

cyclonev_lcell_comb \sr[14]~10 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[14]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[14]~10 .extended_lut = "off";
defparam \sr[14]~10 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \sr[14]~10 .shared_arith = "off";

cyclonev_lcell_comb \sr~11 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_3),
	.datad(!break_readreg_1),
	.datae(!MonDReg_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~11 .extended_lut = "off";
defparam \sr~11 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~11 .shared_arith = "off";

cyclonev_lcell_comb \sr~12 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_4),
	.datad(!break_readreg_2),
	.datae(!MonDReg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~12 .extended_lut = "off";
defparam \sr~12 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~12 .shared_arith = "off";

cyclonev_lcell_comb \sr~13 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_5),
	.datad(!break_readreg_3),
	.datae(!MonDReg_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~13 .extended_lut = "off";
defparam \sr~13 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~13 .shared_arith = "off";

cyclonev_lcell_comb \sr~20 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_18),
	.datad(!break_readreg_16),
	.datae(!MonDReg_16),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~20 .extended_lut = "off";
defparam \sr~20 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~20 .shared_arith = "off";

cyclonev_lcell_comb \sr[29]~21 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!irf_reg_0_2),
	.datae(!irf_reg_1_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[29]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[29]~21 .extended_lut = "off";
defparam \sr[29]~21 .lut_mask = 64'hFFFFFBFFFFFFFBFF;
defparam \sr[29]~21 .shared_arith = "off";

cyclonev_lcell_comb \sr[29]~19 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(!irf_reg_0_2),
	.dataf(!irf_reg_1_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[29]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[29]~19 .extended_lut = "off";
defparam \sr[29]~19 .lut_mask = 64'hFFFFFFFFFFFFDFFF;
defparam \sr[29]~19 .shared_arith = "off";

cyclonev_lcell_comb \sr~22 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_26),
	.datad(!break_readreg_24),
	.datae(!MonDReg_24),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~22 .extended_lut = "off";
defparam \sr~22 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~22 .shared_arith = "off";

cyclonev_lcell_comb \sr~23 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_6),
	.datad(!break_readreg_4),
	.datae(!MonDReg_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~23 .extended_lut = "off";
defparam \sr~23 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~23 .shared_arith = "off";

cyclonev_lcell_comb \sr~24 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_27),
	.datad(!break_readreg_25),
	.datae(!MonDReg_25),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~24 .extended_lut = "off";
defparam \sr~24 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~24 .shared_arith = "off";

cyclonev_lcell_comb \sr~25 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_29),
	.datad(!break_readreg_27),
	.datae(!MonDReg_27),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~25 .extended_lut = "off";
defparam \sr~25 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~25 .shared_arith = "off";

cyclonev_lcell_comb \sr~26 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_28),
	.datad(!break_readreg_26),
	.datae(!MonDReg_26),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~26 .extended_lut = "off";
defparam \sr~26 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~26 .shared_arith = "off";

cyclonev_lcell_comb \sr~27 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_22),
	.datad(!break_readreg_20),
	.datae(!MonDReg_20),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~27 .extended_lut = "off";
defparam \sr~27 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~27 .shared_arith = "off";

cyclonev_lcell_comb \sr~28 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_21),
	.datad(!break_readreg_19),
	.datae(!MonDReg_19),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~28 .extended_lut = "off";
defparam \sr~28 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~28 .shared_arith = "off";

cyclonev_lcell_comb \sr~29 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_19),
	.datad(!MonDReg_17),
	.datae(!break_readreg_17),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~29 .extended_lut = "off";
defparam \sr~29 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~29 .shared_arith = "off";

cyclonev_lcell_comb \sr~30 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_5),
	.datad(!sr_7),
	.datae(!break_readreg_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~30 .extended_lut = "off";
defparam \sr~30 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~30 .shared_arith = "off";

cyclonev_lcell_comb \sr~31 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_30),
	.datad(!break_readreg_28),
	.datae(!MonDReg_28),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~31 .extended_lut = "off";
defparam \sr~31 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~31 .shared_arith = "off";

cyclonev_lcell_comb \sr~32 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_31),
	.datad(!break_readreg_29),
	.datae(!MonDReg_29),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~32 .extended_lut = "off";
defparam \sr~32 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~32 .shared_arith = "off";

cyclonev_lcell_comb \sr~37 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_33),
	.datad(!break_readreg_31),
	.datae(!MonDReg_31),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~37 .extended_lut = "off";
defparam \sr~37 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~37 .shared_arith = "off";

cyclonev_lcell_comb \sr~39 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_21),
	.datad(!sr_23),
	.datae(!break_readreg_21),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~39 .extended_lut = "off";
defparam \sr~39 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~39 .shared_arith = "off";

cyclonev_lcell_comb \sr~40 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_20),
	.datad(!MonDReg_18),
	.datae(!break_readreg_18),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~40 .extended_lut = "off";
defparam \sr~40 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~40 .shared_arith = "off";

cyclonev_lcell_comb \sr~43 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_22),
	.datad(!sr_24),
	.datae(!break_readreg_22),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~43 .extended_lut = "off";
defparam \sr~43 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~43 .shared_arith = "off";

cyclonev_lcell_comb \sr~44 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_17),
	.datad(!MonDReg_15),
	.datae(!break_readreg_15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~44 .extended_lut = "off";
defparam \sr~44 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~44 .shared_arith = "off";

cyclonev_lcell_comb \sr~45 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_25),
	.datad(!MonDReg_23),
	.datae(!break_readreg_23),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~45 .extended_lut = "off";
defparam \sr~45 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~45 .shared_arith = "off";

cyclonev_lcell_comb \sr~46 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_7),
	.datad(!sr_9),
	.datae(!break_readreg_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~46 .extended_lut = "off";
defparam \sr~46 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~46 .shared_arith = "off";

cyclonev_lcell_comb \sr~47 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_13),
	.datad(!sr_15),
	.datae(!break_readreg_13),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~47 .extended_lut = "off";
defparam \sr~47 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~47 .shared_arith = "off";

cyclonev_lcell_comb \sr~50 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_10),
	.datad(!sr_12),
	.datae(!break_readreg_10),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~50 .extended_lut = "off";
defparam \sr~50 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~50 .shared_arith = "off";

cyclonev_lcell_comb \sr~51 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_12),
	.datad(!sr_14),
	.datae(!break_readreg_12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~51 .extended_lut = "off";
defparam \sr~51 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~51 .shared_arith = "off";

cyclonev_lcell_comb \sr~52 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_11),
	.datad(!sr_13),
	.datae(!break_readreg_11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~52 .extended_lut = "off";
defparam \sr~52 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~52 .shared_arith = "off";

cyclonev_lcell_comb \sr~53 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_8),
	.datad(!sr_10),
	.datae(!break_readreg_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~53 .extended_lut = "off";
defparam \sr~53 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~53 .shared_arith = "off";

cyclonev_lcell_comb \sr~54 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_9),
	.datad(!sr_11),
	.datae(!break_readreg_9),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~54 .extended_lut = "off";
defparam \sr~54 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~54 .shared_arith = "off";

cyclonev_lcell_comb \sr~5 (
	.dataa(!sr_0),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~5 .extended_lut = "off";
defparam \sr~5 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \sr~5 .shared_arith = "off";

cyclonev_lcell_comb \sr~6 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(!\the_altera_std_synchronizer2|dreg[0]~q ),
	.datae(!irf_reg_0_2),
	.dataf(!irf_reg_1_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~6 .extended_lut = "off";
defparam \sr~6 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \sr~6 .shared_arith = "off";

dffeas \DRsize.000 (
	.clk(altera_internal_jtag),
	.d(vcc),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.000~q ),
	.prn(vcc));
defparam \DRsize.000 .is_wysiwyg = "true";
defparam \DRsize.000 .power_up = "low";

cyclonev_lcell_comb \sr~7 (
	.dataa(!virtual_state_sdr),
	.datab(!\sr~5_combout ),
	.datac(!\sr~6_combout ),
	.datad(!sr_1),
	.datae(!\DRsize.000~q ),
	.dataf(!altera_internal_jtag1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~7 .extended_lut = "off";
defparam \sr~7 .lut_mask = 64'h7FFFBFFFFFFFFFFF;
defparam \sr~7 .shared_arith = "off";

cyclonev_lcell_comb \sr~14 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!sr_37),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~14 .extended_lut = "off";
defparam \sr~14 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \sr~14 .shared_arith = "off";

cyclonev_lcell_comb \sr[37]~15 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(!irf_reg_0_2),
	.dataf(!irf_reg_1_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[37]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[37]~15 .extended_lut = "off";
defparam \sr[37]~15 .lut_mask = 64'hDFFFFFFFFFFFDFFF;
defparam \sr[37]~15 .shared_arith = "off";

cyclonev_lcell_comb \sr~16 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!altera_internal_jtag1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~16 .extended_lut = "off";
defparam \sr~16 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \sr~16 .shared_arith = "off";

cyclonev_lcell_comb \Mux37~0 (
	.dataa(!irf_reg_0_2),
	.datab(!irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux37~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux37~0 .extended_lut = "off";
defparam \Mux37~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Mux37~0 .shared_arith = "off";

dffeas \DRsize.100 (
	.clk(altera_internal_jtag),
	.d(\Mux37~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.100~q ),
	.prn(vcc));
defparam \DRsize.100 .is_wysiwyg = "true";
defparam \DRsize.100 .power_up = "low";

cyclonev_lcell_comb \sr~56 (
	.dataa(!virtual_state_cdr),
	.datab(!sr_35),
	.datac(!irf_reg_0_2),
	.datad(!irf_reg_1_2),
	.datae(!\the_altera_std_synchronizer1|dreg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~56 .extended_lut = "off";
defparam \sr~56 .lut_mask = 64'hB77BFFFFB77BFFFF;
defparam \sr~56 .shared_arith = "off";

cyclonev_lcell_comb \sr~17 (
	.dataa(!virtual_state_sdr),
	.datab(!altera_internal_jtag1),
	.datac(!sr_36),
	.datad(!\DRsize.100~q ),
	.datae(!\sr~56_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~17 .extended_lut = "off";
defparam \sr~17 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \sr~17 .shared_arith = "off";

cyclonev_lcell_comb \sr~18 (
	.dataa(!virtual_state_sdr),
	.datab(!\Mux37~0_combout ),
	.datac(!sr_35),
	.datad(!monitor_error),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~18 .extended_lut = "off";
defparam \sr~18 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \sr~18 .shared_arith = "off";

cyclonev_lcell_comb \sr[29]~33 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(!irf_reg_0_2),
	.datae(!irf_reg_1_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[29]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[29]~33 .extended_lut = "off";
defparam \sr[29]~33 .lut_mask = 64'hFFFFFFBFFFFFFFBF;
defparam \sr[29]~33 .shared_arith = "off";

cyclonev_lcell_comb \sr~34 (
	.dataa(!irf_reg_1_2),
	.datab(!MonDReg_30),
	.datac(!break_readreg_30),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~34 .extended_lut = "off";
defparam \sr~34 .lut_mask = 64'h2727272727272727;
defparam \sr~34 .shared_arith = "off";

cyclonev_lcell_comb \sr~35 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(!irf_reg_0_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~35 .extended_lut = "off";
defparam \sr~35 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \sr~35 .shared_arith = "off";

cyclonev_lcell_comb \sr~36 (
	.dataa(!virtual_state_sdr),
	.datab(!\sr[29]~33_combout ),
	.datac(!sr_31),
	.datad(!sr_32),
	.datae(!\sr~34_combout ),
	.dataf(!\sr~35_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~36 .extended_lut = "off";
defparam \sr~36 .lut_mask = 64'h8DFFFFFFFFFFFFFF;
defparam \sr~36 .shared_arith = "off";

cyclonev_lcell_comb \sr~38 (
	.dataa(!virtual_state_sdr),
	.datab(!\Mux37~0_combout ),
	.datac(!sr_34),
	.datad(!resetlatch),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~38 .extended_lut = "off";
defparam \sr~38 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \sr~38 .shared_arith = "off";

cyclonev_lcell_comb \sr~41 (
	.dataa(!irf_reg_1_2),
	.datab(!MonDReg_6),
	.datac(!break_readreg_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~41 .extended_lut = "off";
defparam \sr~41 .lut_mask = 64'h2727272727272727;
defparam \sr~41 .shared_arith = "off";

cyclonev_lcell_comb \sr~42 (
	.dataa(!virtual_state_sdr),
	.datab(!virtual_state_cdr),
	.datac(!irf_reg_0_2),
	.datad(!sr_7),
	.datae(!sr_8),
	.dataf(!\sr~41_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~42 .extended_lut = "off";
defparam \sr~42 .lut_mask = 64'hF6FFFFFFFFFFFFFF;
defparam \sr~42 .shared_arith = "off";

cyclonev_lcell_comb \sr[29]~55 (
	.dataa(!irf_reg_0_2),
	.datab(!irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[29]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[29]~55 .extended_lut = "off";
defparam \sr[29]~55 .lut_mask = 64'h7777777777777777;
defparam \sr[29]~55 .shared_arith = "off";

dffeas \DRsize.010 (
	.clk(altera_internal_jtag),
	.d(\sr[29]~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.010~q ),
	.prn(vcc));
defparam \DRsize.010 .is_wysiwyg = "true";
defparam \DRsize.010 .power_up = "low";

cyclonev_lcell_comb \sr~48 (
	.dataa(!virtual_state_cdr),
	.datab(!irf_reg_0_2),
	.datac(!irf_reg_1_2),
	.datad(!MonDReg_14),
	.datae(!sr_15),
	.dataf(!break_readreg_14),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~48 .extended_lut = "off";
defparam \sr~48 .lut_mask = 64'hDEFFFFFFFFFFFFFF;
defparam \sr~48 .shared_arith = "off";

cyclonev_lcell_comb \sr~49 (
	.dataa(!virtual_state_sdr),
	.datab(!altera_internal_jtag1),
	.datac(!sr_16),
	.datad(!\DRsize.010~q ),
	.datae(!\sr~48_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~49 .extended_lut = "off";
defparam \sr~49 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \sr~49 .shared_arith = "off";

endmodule

module niosLab2_altera_std_synchronizer_2 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosLab2_altera_std_synchronizer_3 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosLab2_sld_virtual_jtag_basic_1 (
	virtual_state_sdr,
	virtual_state_uir1,
	virtual_state_cdr1,
	virtual_state_udr,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3)/* synthesis synthesis_greybox=1 */;
output 	virtual_state_sdr;
output 	virtual_state_uir1;
output 	virtual_state_cdr1;
output 	virtual_state_udr;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \virtual_state_sdr~0 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_sdr),
	.sumout(),
	.cout(),
	.shareout());
defparam \virtual_state_sdr~0 .extended_lut = "off";
defparam \virtual_state_sdr~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \virtual_state_sdr~0 .shared_arith = "off";

cyclonev_lcell_comb virtual_state_uir(
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_uir1),
	.sumout(),
	.cout(),
	.shareout());
defparam virtual_state_uir.extended_lut = "off";
defparam virtual_state_uir.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam virtual_state_uir.shared_arith = "off";

cyclonev_lcell_comb virtual_state_cdr(
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_cdr1),
	.sumout(),
	.cout(),
	.shareout());
defparam virtual_state_cdr.extended_lut = "off";
defparam virtual_state_cdr.lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam virtual_state_cdr.shared_arith = "off";

cyclonev_lcell_comb \virtual_state_udr~0 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_udr),
	.sumout(),
	.cout(),
	.shareout());
defparam \virtual_state_udr~0 .extended_lut = "off";
defparam \virtual_state_udr~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \virtual_state_udr~0 .shared_arith = "off";

endmodule

module niosLab2_niosLab2_nios2_gen2_0_cpu_nios2_avalon_reg (
	r_sync_rst,
	write,
	address_8,
	address_0,
	address_3,
	address_7,
	address_6,
	address_5,
	address_4,
	address_2,
	address_1,
	debugaccess,
	take_action_ocireg,
	oci_single_step_mode1,
	Equal0,
	oci_ienable_16,
	oci_reg_readdata,
	writedata_3,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	write;
input 	address_8;
input 	address_0;
input 	address_3;
input 	address_7;
input 	address_6;
input 	address_5;
input 	address_4;
input 	address_2;
input 	address_1;
input 	debugaccess;
output 	take_action_ocireg;
output 	oci_single_step_mode1;
output 	Equal0;
output 	oci_ienable_16;
output 	oci_reg_readdata;
input 	writedata_3;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \oci_single_step_mode~0_combout ;
wire \oci_ienable[16]~0_combout ;


cyclonev_lcell_comb \take_action_ocireg~0 (
	.dataa(!write),
	.datab(!address_0),
	.datac(!address_3),
	.datad(!\Equal0~0_combout ),
	.datae(!\Equal0~1_combout ),
	.dataf(!debugaccess),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocireg),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_ocireg~0 .extended_lut = "off";
defparam \take_action_ocireg~0 .lut_mask = 64'hFDFFFFFFFFFFFFFF;
defparam \take_action_ocireg~0 .shared_arith = "off";

dffeas oci_single_step_mode(
	.clk(clk_clk),
	.d(\oci_single_step_mode~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oci_single_step_mode1),
	.prn(vcc));
defparam oci_single_step_mode.is_wysiwyg = "true";
defparam oci_single_step_mode.power_up = "low";

cyclonev_lcell_comb \Equal0~2 (
	.dataa(!address_3),
	.datab(!\Equal0~0_combout ),
	.datac(!\Equal0~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~2 .extended_lut = "off";
defparam \Equal0~2 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \Equal0~2 .shared_arith = "off";

dffeas \oci_ienable[16] (
	.clk(clk_clk),
	.d(\oci_ienable[16]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oci_ienable_16),
	.prn(vcc));
defparam \oci_ienable[16] .is_wysiwyg = "true";
defparam \oci_ienable[16] .power_up = "low";

cyclonev_lcell_comb \oci_reg_readdata~0 (
	.dataa(!address_0),
	.datab(!Equal0),
	.datac(!oci_ienable_16),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(oci_reg_readdata),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_reg_readdata~0 .extended_lut = "off";
defparam \oci_reg_readdata~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \oci_reg_readdata~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!address_8),
	.datab(!address_7),
	.datac(!address_6),
	.datad(!address_5),
	.datae(!address_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!address_2),
	.datab(!address_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \oci_single_step_mode~0 (
	.dataa(!take_action_ocireg),
	.datab(!oci_single_step_mode1),
	.datac(!writedata_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\oci_single_step_mode~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_single_step_mode~0 .extended_lut = "off";
defparam \oci_single_step_mode~0 .lut_mask = 64'h2727272727272727;
defparam \oci_single_step_mode~0 .shared_arith = "off";

cyclonev_lcell_comb \oci_ienable[16]~0 (
	.dataa(!write),
	.datab(!address_0),
	.datac(!Equal0),
	.datad(!debugaccess),
	.datae(!oci_ienable_16),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\oci_ienable[16]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_ienable[16]~0 .extended_lut = "off";
defparam \oci_ienable[16]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \oci_ienable[16]~0 .shared_arith = "off";

endmodule

module niosLab2_niosLab2_nios2_gen2_0_cpu_nios2_oci_break (
	break_readreg_0,
	break_readreg_1,
	break_readreg_2,
	break_readreg_3,
	break_readreg_16,
	break_readreg_24,
	break_readreg_4,
	break_readreg_25,
	break_readreg_27,
	break_readreg_26,
	break_readreg_20,
	break_readreg_19,
	break_readreg_17,
	break_readreg_5,
	break_readreg_28,
	break_readreg_29,
	break_readreg_30,
	break_readreg_31,
	break_readreg_21,
	break_readreg_18,
	break_readreg_6,
	break_readreg_22,
	break_readreg_15,
	break_readreg_23,
	break_readreg_7,
	break_readreg_13,
	break_readreg_14,
	break_readreg_10,
	break_readreg_12,
	break_readreg_11,
	break_readreg_8,
	break_readreg_9,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_1,
	ir_0,
	enable_action_strobe,
	jdo_3,
	jdo_17,
	jdo_25,
	jdo_1,
	jdo_4,
	jdo_26,
	jdo_28,
	jdo_27,
	jdo_21,
	jdo_20,
	jdo_2,
	jdo_5,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_19,
	jdo_18,
	jdo_6,
	jdo_23,
	jdo_16,
	jdo_24,
	jdo_7,
	jdo_22,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_11,
	jdo_13,
	jdo_12,
	jdo_9,
	jdo_10,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	break_readreg_0;
output 	break_readreg_1;
output 	break_readreg_2;
output 	break_readreg_3;
output 	break_readreg_16;
output 	break_readreg_24;
output 	break_readreg_4;
output 	break_readreg_25;
output 	break_readreg_27;
output 	break_readreg_26;
output 	break_readreg_20;
output 	break_readreg_19;
output 	break_readreg_17;
output 	break_readreg_5;
output 	break_readreg_28;
output 	break_readreg_29;
output 	break_readreg_30;
output 	break_readreg_31;
output 	break_readreg_21;
output 	break_readreg_18;
output 	break_readreg_6;
output 	break_readreg_22;
output 	break_readreg_15;
output 	break_readreg_23;
output 	break_readreg_7;
output 	break_readreg_13;
output 	break_readreg_14;
output 	break_readreg_10;
output 	break_readreg_12;
output 	break_readreg_11;
output 	break_readreg_8;
output 	break_readreg_9;
input 	jdo_0;
input 	jdo_36;
input 	jdo_37;
input 	ir_1;
input 	ir_0;
input 	enable_action_strobe;
input 	jdo_3;
input 	jdo_17;
input 	jdo_25;
input 	jdo_1;
input 	jdo_4;
input 	jdo_26;
input 	jdo_28;
input 	jdo_27;
input 	jdo_21;
input 	jdo_20;
input 	jdo_2;
input 	jdo_5;
input 	jdo_29;
input 	jdo_30;
input 	jdo_31;
input 	jdo_19;
input 	jdo_18;
input 	jdo_6;
input 	jdo_23;
input 	jdo_16;
input 	jdo_24;
input 	jdo_7;
input 	jdo_22;
input 	jdo_14;
input 	jdo_15;
input 	jdo_8;
input 	jdo_11;
input 	jdo_13;
input 	jdo_12;
input 	jdo_9;
input 	jdo_10;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \break_readreg[13]~0_combout ;
wire \break_readreg[13]~1_combout ;


dffeas \break_readreg[0] (
	.clk(clk_clk),
	.d(jdo_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_0),
	.prn(vcc));
defparam \break_readreg[0] .is_wysiwyg = "true";
defparam \break_readreg[0] .power_up = "low";

dffeas \break_readreg[1] (
	.clk(clk_clk),
	.d(jdo_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_1),
	.prn(vcc));
defparam \break_readreg[1] .is_wysiwyg = "true";
defparam \break_readreg[1] .power_up = "low";

dffeas \break_readreg[2] (
	.clk(clk_clk),
	.d(jdo_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_2),
	.prn(vcc));
defparam \break_readreg[2] .is_wysiwyg = "true";
defparam \break_readreg[2] .power_up = "low";

dffeas \break_readreg[3] (
	.clk(clk_clk),
	.d(jdo_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_3),
	.prn(vcc));
defparam \break_readreg[3] .is_wysiwyg = "true";
defparam \break_readreg[3] .power_up = "low";

dffeas \break_readreg[16] (
	.clk(clk_clk),
	.d(jdo_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_16),
	.prn(vcc));
defparam \break_readreg[16] .is_wysiwyg = "true";
defparam \break_readreg[16] .power_up = "low";

dffeas \break_readreg[24] (
	.clk(clk_clk),
	.d(jdo_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_24),
	.prn(vcc));
defparam \break_readreg[24] .is_wysiwyg = "true";
defparam \break_readreg[24] .power_up = "low";

dffeas \break_readreg[4] (
	.clk(clk_clk),
	.d(jdo_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_4),
	.prn(vcc));
defparam \break_readreg[4] .is_wysiwyg = "true";
defparam \break_readreg[4] .power_up = "low";

dffeas \break_readreg[25] (
	.clk(clk_clk),
	.d(jdo_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_25),
	.prn(vcc));
defparam \break_readreg[25] .is_wysiwyg = "true";
defparam \break_readreg[25] .power_up = "low";

dffeas \break_readreg[27] (
	.clk(clk_clk),
	.d(jdo_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_27),
	.prn(vcc));
defparam \break_readreg[27] .is_wysiwyg = "true";
defparam \break_readreg[27] .power_up = "low";

dffeas \break_readreg[26] (
	.clk(clk_clk),
	.d(jdo_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_26),
	.prn(vcc));
defparam \break_readreg[26] .is_wysiwyg = "true";
defparam \break_readreg[26] .power_up = "low";

dffeas \break_readreg[20] (
	.clk(clk_clk),
	.d(jdo_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_20),
	.prn(vcc));
defparam \break_readreg[20] .is_wysiwyg = "true";
defparam \break_readreg[20] .power_up = "low";

dffeas \break_readreg[19] (
	.clk(clk_clk),
	.d(jdo_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_19),
	.prn(vcc));
defparam \break_readreg[19] .is_wysiwyg = "true";
defparam \break_readreg[19] .power_up = "low";

dffeas \break_readreg[17] (
	.clk(clk_clk),
	.d(jdo_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_17),
	.prn(vcc));
defparam \break_readreg[17] .is_wysiwyg = "true";
defparam \break_readreg[17] .power_up = "low";

dffeas \break_readreg[5] (
	.clk(clk_clk),
	.d(jdo_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_5),
	.prn(vcc));
defparam \break_readreg[5] .is_wysiwyg = "true";
defparam \break_readreg[5] .power_up = "low";

dffeas \break_readreg[28] (
	.clk(clk_clk),
	.d(jdo_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_28),
	.prn(vcc));
defparam \break_readreg[28] .is_wysiwyg = "true";
defparam \break_readreg[28] .power_up = "low";

dffeas \break_readreg[29] (
	.clk(clk_clk),
	.d(jdo_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_29),
	.prn(vcc));
defparam \break_readreg[29] .is_wysiwyg = "true";
defparam \break_readreg[29] .power_up = "low";

dffeas \break_readreg[30] (
	.clk(clk_clk),
	.d(jdo_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_30),
	.prn(vcc));
defparam \break_readreg[30] .is_wysiwyg = "true";
defparam \break_readreg[30] .power_up = "low";

dffeas \break_readreg[31] (
	.clk(clk_clk),
	.d(jdo_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_31),
	.prn(vcc));
defparam \break_readreg[31] .is_wysiwyg = "true";
defparam \break_readreg[31] .power_up = "low";

dffeas \break_readreg[21] (
	.clk(clk_clk),
	.d(jdo_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_21),
	.prn(vcc));
defparam \break_readreg[21] .is_wysiwyg = "true";
defparam \break_readreg[21] .power_up = "low";

dffeas \break_readreg[18] (
	.clk(clk_clk),
	.d(jdo_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_18),
	.prn(vcc));
defparam \break_readreg[18] .is_wysiwyg = "true";
defparam \break_readreg[18] .power_up = "low";

dffeas \break_readreg[6] (
	.clk(clk_clk),
	.d(jdo_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_6),
	.prn(vcc));
defparam \break_readreg[6] .is_wysiwyg = "true";
defparam \break_readreg[6] .power_up = "low";

dffeas \break_readreg[22] (
	.clk(clk_clk),
	.d(jdo_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_22),
	.prn(vcc));
defparam \break_readreg[22] .is_wysiwyg = "true";
defparam \break_readreg[22] .power_up = "low";

dffeas \break_readreg[15] (
	.clk(clk_clk),
	.d(jdo_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_15),
	.prn(vcc));
defparam \break_readreg[15] .is_wysiwyg = "true";
defparam \break_readreg[15] .power_up = "low";

dffeas \break_readreg[23] (
	.clk(clk_clk),
	.d(jdo_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_23),
	.prn(vcc));
defparam \break_readreg[23] .is_wysiwyg = "true";
defparam \break_readreg[23] .power_up = "low";

dffeas \break_readreg[7] (
	.clk(clk_clk),
	.d(jdo_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_7),
	.prn(vcc));
defparam \break_readreg[7] .is_wysiwyg = "true";
defparam \break_readreg[7] .power_up = "low";

dffeas \break_readreg[13] (
	.clk(clk_clk),
	.d(jdo_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_13),
	.prn(vcc));
defparam \break_readreg[13] .is_wysiwyg = "true";
defparam \break_readreg[13] .power_up = "low";

dffeas \break_readreg[14] (
	.clk(clk_clk),
	.d(jdo_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_14),
	.prn(vcc));
defparam \break_readreg[14] .is_wysiwyg = "true";
defparam \break_readreg[14] .power_up = "low";

dffeas \break_readreg[10] (
	.clk(clk_clk),
	.d(jdo_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_10),
	.prn(vcc));
defparam \break_readreg[10] .is_wysiwyg = "true";
defparam \break_readreg[10] .power_up = "low";

dffeas \break_readreg[12] (
	.clk(clk_clk),
	.d(jdo_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_12),
	.prn(vcc));
defparam \break_readreg[12] .is_wysiwyg = "true";
defparam \break_readreg[12] .power_up = "low";

dffeas \break_readreg[11] (
	.clk(clk_clk),
	.d(jdo_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_11),
	.prn(vcc));
defparam \break_readreg[11] .is_wysiwyg = "true";
defparam \break_readreg[11] .power_up = "low";

dffeas \break_readreg[8] (
	.clk(clk_clk),
	.d(jdo_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_8),
	.prn(vcc));
defparam \break_readreg[8] .is_wysiwyg = "true";
defparam \break_readreg[8] .power_up = "low";

dffeas \break_readreg[9] (
	.clk(clk_clk),
	.d(jdo_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[13]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[13]~0_combout ),
	.q(break_readreg_9),
	.prn(vcc));
defparam \break_readreg[9] .is_wysiwyg = "true";
defparam \break_readreg[9] .power_up = "low";

cyclonev_lcell_comb \break_readreg[13]~0 (
	.dataa(!ir_1),
	.datab(!ir_0),
	.datac(!enable_action_strobe),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\break_readreg[13]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \break_readreg[13]~0 .extended_lut = "off";
defparam \break_readreg[13]~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \break_readreg[13]~0 .shared_arith = "off";

cyclonev_lcell_comb \break_readreg[13]~1 (
	.dataa(!jdo_36),
	.datab(!jdo_37),
	.datac(!\break_readreg[13]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\break_readreg[13]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \break_readreg[13]~1 .extended_lut = "off";
defparam \break_readreg[13]~1 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \break_readreg[13]~1 .shared_arith = "off";

endmodule

module niosLab2_niosLab2_nios2_gen2_0_cpu_nios2_oci_debug (
	r_sync_rst,
	monitor_ready1,
	jtag_break1,
	jdo_34,
	take_action_ocimem_a,
	take_action_ocimem_a1,
	jdo_25,
	writedata_0,
	take_action_ocireg,
	jdo_21,
	jdo_20,
	writedata_1,
	monitor_error1,
	jdo_19,
	jdo_18,
	monitor_go1,
	jdo_23,
	jdo_24,
	resetlatch1,
	state_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	monitor_ready1;
output 	jtag_break1;
input 	jdo_34;
input 	take_action_ocimem_a;
input 	take_action_ocimem_a1;
input 	jdo_25;
input 	writedata_0;
input 	take_action_ocireg;
input 	jdo_21;
input 	jdo_20;
input 	writedata_1;
output 	monitor_error1;
input 	jdo_19;
input 	jdo_18;
output 	monitor_go1;
input 	jdo_23;
input 	jdo_24;
output 	resetlatch1;
input 	state_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer|dreg[0]~q ;
wire \monitor_ready~0_combout ;
wire \break_on_reset~0_combout ;
wire \break_on_reset~q ;
wire \jtag_break~0_combout ;
wire \monitor_error~0_combout ;
wire \monitor_go~0_combout ;
wire \resetlatch~0_combout ;


niosLab2_altera_std_synchronizer_4 the_altera_std_synchronizer(
	.din(r_sync_rst),
	.dreg_0(\the_altera_std_synchronizer|dreg[0]~q ),
	.clk(clk_clk));

dffeas monitor_ready(
	.clk(clk_clk),
	.d(\monitor_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_ready1),
	.prn(vcc));
defparam monitor_ready.is_wysiwyg = "true";
defparam monitor_ready.power_up = "low";

dffeas jtag_break(
	.clk(clk_clk),
	.d(\jtag_break~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(jtag_break1),
	.prn(vcc));
defparam jtag_break.is_wysiwyg = "true";
defparam jtag_break.power_up = "low";

dffeas monitor_error(
	.clk(clk_clk),
	.d(\monitor_error~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_error1),
	.prn(vcc));
defparam monitor_error.is_wysiwyg = "true";
defparam monitor_error.power_up = "low";

dffeas monitor_go(
	.clk(clk_clk),
	.d(\monitor_go~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_go1),
	.prn(vcc));
defparam monitor_go.is_wysiwyg = "true";
defparam monitor_go.power_up = "low";

dffeas resetlatch(
	.clk(clk_clk),
	.d(\resetlatch~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(resetlatch1),
	.prn(vcc));
defparam resetlatch.is_wysiwyg = "true";
defparam resetlatch.power_up = "low";

cyclonev_lcell_comb \monitor_ready~0 (
	.dataa(!monitor_ready1),
	.datab(!take_action_ocimem_a1),
	.datac(!jdo_25),
	.datad(!writedata_0),
	.datae(!take_action_ocireg),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\monitor_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \monitor_ready~0 .extended_lut = "off";
defparam \monitor_ready~0 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \monitor_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \break_on_reset~0 (
	.dataa(!take_action_ocimem_a1),
	.datab(!\break_on_reset~q ),
	.datac(!jdo_19),
	.datad(!jdo_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\break_on_reset~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \break_on_reset~0 .extended_lut = "off";
defparam \break_on_reset~0 .lut_mask = 64'hBF1FBF1FBF1FBF1F;
defparam \break_on_reset~0 .shared_arith = "off";

dffeas break_on_reset(
	.clk(clk_clk),
	.d(\break_on_reset~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\break_on_reset~q ),
	.prn(vcc));
defparam break_on_reset.is_wysiwyg = "true";
defparam break_on_reset.power_up = "low";

cyclonev_lcell_comb \jtag_break~0 (
	.dataa(!jtag_break1),
	.datab(!take_action_ocimem_a1),
	.datac(!jdo_21),
	.datad(!jdo_20),
	.datae(!\break_on_reset~q ),
	.dataf(!\the_altera_std_synchronizer|dreg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_break~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_break~0 .extended_lut = "off";
defparam \jtag_break~0 .lut_mask = 64'hFF7FFFFFFFDFFFFF;
defparam \jtag_break~0 .shared_arith = "off";

cyclonev_lcell_comb \monitor_error~0 (
	.dataa(!take_action_ocimem_a1),
	.datab(!jdo_25),
	.datac(!take_action_ocireg),
	.datad(!writedata_1),
	.datae(!monitor_error1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\monitor_error~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \monitor_error~0 .extended_lut = "off";
defparam \monitor_error~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \monitor_error~0 .shared_arith = "off";

cyclonev_lcell_comb \monitor_go~0 (
	.dataa(!take_action_ocimem_a),
	.datab(!jdo_34),
	.datac(!monitor_go1),
	.datad(!jdo_23),
	.datae(!state_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\monitor_go~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \monitor_go~0 .extended_lut = "off";
defparam \monitor_go~0 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \monitor_go~0 .shared_arith = "off";

cyclonev_lcell_comb \resetlatch~0 (
	.dataa(!take_action_ocimem_a1),
	.datab(!\the_altera_std_synchronizer|dreg[0]~q ),
	.datac(!jdo_24),
	.datad(!resetlatch1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\resetlatch~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \resetlatch~0 .extended_lut = "off";
defparam \resetlatch~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \resetlatch~0 .shared_arith = "off";

endmodule

module niosLab2_altera_std_synchronizer_4 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module niosLab2_niosLab2_nios2_gen2_0_cpu_nios2_ocimem (
	MonDReg_1,
	q_a_0,
	MonDReg_2,
	q_a_1,
	MonDReg_3,
	q_a_2,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_11,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_15,
	q_a_16,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_8,
	q_a_10,
	q_a_17,
	q_a_9,
	q_a_18,
	q_a_19,
	q_a_20,
	q_a_21,
	q_a_6,
	MonDReg_16,
	q_a_7,
	MonDReg_24,
	MonDReg_25,
	MonDReg_27,
	MonDReg_26,
	MonDReg_22,
	MonDReg_20,
	MonDReg_19,
	MonDReg_23,
	MonDReg_11,
	MonDReg_13,
	MonDReg_14,
	q_a_27,
	q_a_28,
	q_a_29,
	q_a_30,
	q_a_31,
	MonDReg_10,
	MonDReg_17,
	MonDReg_9,
	MonDReg_21,
	MonDReg_6,
	MonDReg_7,
	MonDReg_28,
	MonDReg_30,
	MonDReg_31,
	waitrequest1,
	MonDReg_0,
	write,
	address_8,
	read,
	ir_1,
	ir_0,
	enable_action_strobe,
	jdo_35,
	take_action_ocimem_b,
	jdo_3,
	take_action_ocimem_a,
	jdo_34,
	jdo_17,
	take_action_ocimem_a1,
	take_action_ocimem_a2,
	jdo_25,
	writedata_0,
	address_0,
	address_3,
	address_7,
	address_6,
	address_5,
	address_4,
	address_2,
	address_1,
	debugaccess,
	jdo_4,
	r_early_rst,
	byteenable_0,
	jdo_26,
	jdo_28,
	jdo_27,
	jdo_21,
	jdo_20,
	jdo_5,
	writedata_1,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	jdo_19,
	jdo_18,
	writedata_3,
	MonDReg_4,
	jdo_6,
	writedata_2,
	writedata_22,
	byteenable_2,
	writedata_23,
	writedata_24,
	byteenable_3,
	writedata_25,
	writedata_26,
	writedata_11,
	byteenable_1,
	MonDReg_12,
	writedata_12,
	writedata_13,
	writedata_14,
	MonDReg_15,
	writedata_15,
	writedata_16,
	jdo_23,
	writedata_4,
	MonDReg_5,
	writedata_5,
	MonDReg_8,
	writedata_8,
	writedata_10,
	writedata_17,
	writedata_9,
	MonDReg_18,
	writedata_18,
	writedata_19,
	writedata_20,
	writedata_21,
	writedata_6,
	jdo_16,
	writedata_7,
	jdo_24,
	jdo_7,
	MonDReg_29,
	jdo_22,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_11,
	writedata_27,
	writedata_28,
	writedata_29,
	writedata_30,
	writedata_31,
	jdo_13,
	jdo_12,
	jdo_9,
	jdo_10,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	MonDReg_1;
output 	q_a_0;
output 	MonDReg_2;
output 	q_a_1;
output 	MonDReg_3;
output 	q_a_2;
output 	q_a_22;
output 	q_a_23;
output 	q_a_24;
output 	q_a_25;
output 	q_a_26;
output 	q_a_11;
output 	q_a_12;
output 	q_a_13;
output 	q_a_14;
output 	q_a_15;
output 	q_a_16;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_8;
output 	q_a_10;
output 	q_a_17;
output 	q_a_9;
output 	q_a_18;
output 	q_a_19;
output 	q_a_20;
output 	q_a_21;
output 	q_a_6;
output 	MonDReg_16;
output 	q_a_7;
output 	MonDReg_24;
output 	MonDReg_25;
output 	MonDReg_27;
output 	MonDReg_26;
output 	MonDReg_22;
output 	MonDReg_20;
output 	MonDReg_19;
output 	MonDReg_23;
output 	MonDReg_11;
output 	MonDReg_13;
output 	MonDReg_14;
output 	q_a_27;
output 	q_a_28;
output 	q_a_29;
output 	q_a_30;
output 	q_a_31;
output 	MonDReg_10;
output 	MonDReg_17;
output 	MonDReg_9;
output 	MonDReg_21;
output 	MonDReg_6;
output 	MonDReg_7;
output 	MonDReg_28;
output 	MonDReg_30;
output 	MonDReg_31;
output 	waitrequest1;
output 	MonDReg_0;
input 	write;
input 	address_8;
input 	read;
input 	ir_1;
input 	ir_0;
input 	enable_action_strobe;
input 	jdo_35;
input 	take_action_ocimem_b;
input 	jdo_3;
input 	take_action_ocimem_a;
input 	jdo_34;
input 	jdo_17;
input 	take_action_ocimem_a1;
input 	take_action_ocimem_a2;
input 	jdo_25;
input 	writedata_0;
input 	address_0;
input 	address_3;
input 	address_7;
input 	address_6;
input 	address_5;
input 	address_4;
input 	address_2;
input 	address_1;
input 	debugaccess;
input 	jdo_4;
input 	r_early_rst;
input 	byteenable_0;
input 	jdo_26;
input 	jdo_28;
input 	jdo_27;
input 	jdo_21;
input 	jdo_20;
input 	jdo_5;
input 	writedata_1;
input 	jdo_29;
input 	jdo_30;
input 	jdo_31;
input 	jdo_32;
input 	jdo_33;
input 	jdo_19;
input 	jdo_18;
input 	writedata_3;
output 	MonDReg_4;
input 	jdo_6;
input 	writedata_2;
input 	writedata_22;
input 	byteenable_2;
input 	writedata_23;
input 	writedata_24;
input 	byteenable_3;
input 	writedata_25;
input 	writedata_26;
input 	writedata_11;
input 	byteenable_1;
output 	MonDReg_12;
input 	writedata_12;
input 	writedata_13;
input 	writedata_14;
output 	MonDReg_15;
input 	writedata_15;
input 	writedata_16;
input 	jdo_23;
input 	writedata_4;
output 	MonDReg_5;
input 	writedata_5;
output 	MonDReg_8;
input 	writedata_8;
input 	writedata_10;
input 	writedata_17;
input 	writedata_9;
output 	MonDReg_18;
input 	writedata_18;
input 	writedata_19;
input 	writedata_20;
input 	writedata_21;
input 	writedata_6;
input 	jdo_16;
input 	writedata_7;
input 	jdo_24;
input 	jdo_7;
output 	MonDReg_29;
input 	jdo_22;
input 	jdo_14;
input 	jdo_15;
input 	jdo_8;
input 	jdo_11;
input 	writedata_27;
input 	writedata_28;
input 	writedata_29;
input 	writedata_30;
input 	writedata_31;
input 	jdo_13;
input 	jdo_12;
input 	jdo_9;
input 	jdo_10;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \jtag_ram_wr~q ;
wire \ociram_wr_en~0_combout ;
wire \ociram_reset_req~combout ;
wire \ociram_wr_data[0]~0_combout ;
wire \ociram_addr[0]~0_combout ;
wire \ociram_addr[1]~1_combout ;
wire \ociram_addr[2]~2_combout ;
wire \ociram_addr[3]~3_combout ;
wire \ociram_addr[4]~4_combout ;
wire \ociram_addr[5]~5_combout ;
wire \ociram_addr[6]~6_combout ;
wire \ociram_addr[7]~7_combout ;
wire \ociram_byteenable[0]~0_combout ;
wire \ociram_wr_data[1]~1_combout ;
wire \jtag_ram_wr~0_combout ;
wire \ociram_wr_data[2]~2_combout ;
wire \ociram_wr_data[22]~3_combout ;
wire \ociram_byteenable[2]~1_combout ;
wire \ociram_wr_data[23]~4_combout ;
wire \ociram_wr_data[24]~5_combout ;
wire \ociram_byteenable[3]~2_combout ;
wire \ociram_wr_data[25]~6_combout ;
wire \ociram_wr_data[26]~7_combout ;
wire \ociram_wr_data[11]~8_combout ;
wire \ociram_byteenable[1]~3_combout ;
wire \ociram_wr_data[12]~9_combout ;
wire \ociram_wr_data[13]~10_combout ;
wire \ociram_wr_data[14]~11_combout ;
wire \ociram_wr_data[15]~12_combout ;
wire \ociram_wr_data[16]~13_combout ;
wire \ociram_wr_data[3]~14_combout ;
wire \ociram_wr_data[4]~15_combout ;
wire \ociram_wr_data[5]~16_combout ;
wire \ociram_wr_data[8]~17_combout ;
wire \ociram_wr_data[10]~18_combout ;
wire \ociram_wr_data[17]~19_combout ;
wire \ociram_wr_data[9]~20_combout ;
wire \ociram_wr_data[18]~21_combout ;
wire \ociram_wr_data[19]~22_combout ;
wire \ociram_wr_data[20]~23_combout ;
wire \ociram_wr_data[21]~24_combout ;
wire \ociram_wr_data[6]~25_combout ;
wire \ociram_wr_data[7]~26_combout ;
wire \ociram_wr_data[27]~27_combout ;
wire \ociram_wr_data[28]~28_combout ;
wire \ociram_wr_data[29]~29_combout ;
wire \ociram_wr_data[30]~30_combout ;
wire \ociram_wr_data[31]~31_combout ;
wire \Add0~1_wirecell_combout ;
wire \MonAReg[10]~q ;
wire \Add0~5_sumout ;
wire \MonAReg[2]~q ;
wire \Add0~6 ;
wire \Add0~13_sumout ;
wire \MonAReg[3]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \MonAReg[4]~q ;
wire \Add0~10 ;
wire \Add0~21_sumout ;
wire \MonAReg[5]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \MonAReg[6]~q ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \MonAReg[7]~q ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \MonAReg[8]~q ;
wire \Add0~34 ;
wire \Add0~17_sumout ;
wire \MonAReg[9]~q ;
wire \Add0~18 ;
wire \Add0~1_sumout ;
wire \jtag_ram_rd~0_combout ;
wire \jtag_ram_rd~q ;
wire \jtag_ram_rd_d1~q ;
wire \MonDReg[11]~3_combout ;
wire \jtag_rd~q ;
wire \jtag_rd_d1~q ;
wire \MonDReg[0]~2_combout ;
wire \jtag_ram_access~0_combout ;
wire \jtag_ram_access~q ;
wire \waitrequest~0_combout ;
wire \avalon_ociram_readdata_ready~0_combout ;
wire \avalon_ociram_readdata_ready~q ;
wire \waitrequest~1_combout ;
wire \MonDReg~0_combout ;
wire \MonDReg~1_combout ;
wire \MonDReg~4_combout ;
wire \MonDReg~5_combout ;
wire \MonDReg[15]~20_combout ;
wire \MonDReg[15]~6_combout ;
wire \MonDReg~16_combout ;
wire \MonDReg[8]~7_combout ;
wire \MonDReg~12_combout ;
wire \MonDReg~8_combout ;


niosLab2_niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module niosLab2_nios2_gen2_0_cpu_ociram_sp_ram(
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_22(q_a_22),
	.q_a_23(q_a_23),
	.q_a_24(q_a_24),
	.q_a_25(q_a_25),
	.q_a_26(q_a_26),
	.q_a_11(q_a_11),
	.q_a_12(q_a_12),
	.q_a_13(q_a_13),
	.q_a_14(q_a_14),
	.q_a_15(q_a_15),
	.q_a_16(q_a_16),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_8(q_a_8),
	.q_a_10(q_a_10),
	.q_a_17(q_a_17),
	.q_a_9(q_a_9),
	.q_a_18(q_a_18),
	.q_a_19(q_a_19),
	.q_a_20(q_a_20),
	.q_a_21(q_a_21),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.q_a_27(q_a_27),
	.q_a_28(q_a_28),
	.q_a_29(q_a_29),
	.q_a_30(q_a_30),
	.q_a_31(q_a_31),
	.ociram_wr_en(\ociram_wr_en~0_combout ),
	.ociram_reset_req(\ociram_reset_req~combout ),
	.ociram_wr_data_0(\ociram_wr_data[0]~0_combout ),
	.ociram_addr_0(\ociram_addr[0]~0_combout ),
	.ociram_addr_1(\ociram_addr[1]~1_combout ),
	.ociram_addr_2(\ociram_addr[2]~2_combout ),
	.ociram_addr_3(\ociram_addr[3]~3_combout ),
	.ociram_addr_4(\ociram_addr[4]~4_combout ),
	.ociram_addr_5(\ociram_addr[5]~5_combout ),
	.ociram_addr_6(\ociram_addr[6]~6_combout ),
	.ociram_addr_7(\ociram_addr[7]~7_combout ),
	.ociram_byteenable_0(\ociram_byteenable[0]~0_combout ),
	.ociram_wr_data_1(\ociram_wr_data[1]~1_combout ),
	.ociram_wr_data_2(\ociram_wr_data[2]~2_combout ),
	.ociram_wr_data_22(\ociram_wr_data[22]~3_combout ),
	.ociram_byteenable_2(\ociram_byteenable[2]~1_combout ),
	.ociram_wr_data_23(\ociram_wr_data[23]~4_combout ),
	.ociram_wr_data_24(\ociram_wr_data[24]~5_combout ),
	.ociram_byteenable_3(\ociram_byteenable[3]~2_combout ),
	.ociram_wr_data_25(\ociram_wr_data[25]~6_combout ),
	.ociram_wr_data_26(\ociram_wr_data[26]~7_combout ),
	.ociram_wr_data_11(\ociram_wr_data[11]~8_combout ),
	.ociram_byteenable_1(\ociram_byteenable[1]~3_combout ),
	.ociram_wr_data_12(\ociram_wr_data[12]~9_combout ),
	.ociram_wr_data_13(\ociram_wr_data[13]~10_combout ),
	.ociram_wr_data_14(\ociram_wr_data[14]~11_combout ),
	.ociram_wr_data_15(\ociram_wr_data[15]~12_combout ),
	.ociram_wr_data_16(\ociram_wr_data[16]~13_combout ),
	.ociram_wr_data_3(\ociram_wr_data[3]~14_combout ),
	.ociram_wr_data_4(\ociram_wr_data[4]~15_combout ),
	.ociram_wr_data_5(\ociram_wr_data[5]~16_combout ),
	.ociram_wr_data_8(\ociram_wr_data[8]~17_combout ),
	.ociram_wr_data_10(\ociram_wr_data[10]~18_combout ),
	.ociram_wr_data_17(\ociram_wr_data[17]~19_combout ),
	.ociram_wr_data_9(\ociram_wr_data[9]~20_combout ),
	.ociram_wr_data_18(\ociram_wr_data[18]~21_combout ),
	.ociram_wr_data_19(\ociram_wr_data[19]~22_combout ),
	.ociram_wr_data_20(\ociram_wr_data[20]~23_combout ),
	.ociram_wr_data_21(\ociram_wr_data[21]~24_combout ),
	.ociram_wr_data_6(\ociram_wr_data[6]~25_combout ),
	.ociram_wr_data_7(\ociram_wr_data[7]~26_combout ),
	.ociram_wr_data_27(\ociram_wr_data[27]~27_combout ),
	.ociram_wr_data_28(\ociram_wr_data[28]~28_combout ),
	.ociram_wr_data_29(\ociram_wr_data[29]~29_combout ),
	.ociram_wr_data_30(\ociram_wr_data[30]~30_combout ),
	.ociram_wr_data_31(\ociram_wr_data[31]~31_combout ),
	.clk_clk(clk_clk));

dffeas jtag_ram_wr(
	.clk(clk_clk),
	.d(\jtag_ram_wr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_wr~q ),
	.prn(vcc));
defparam jtag_ram_wr.is_wysiwyg = "true";
defparam jtag_ram_wr.power_up = "low";

cyclonev_lcell_comb \ociram_wr_en~0 (
	.dataa(!write),
	.datab(!address_8),
	.datac(!\jtag_ram_access~q ),
	.datad(!debugaccess),
	.datae(!\jtag_ram_wr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_en~0 .extended_lut = "off";
defparam \ociram_wr_en~0 .lut_mask = 64'hC5FFFFFFC5FFFFFF;
defparam \ociram_wr_en~0 .shared_arith = "off";

cyclonev_lcell_comb ociram_reset_req(
	.dataa(!\jtag_ram_access~q ),
	.datab(!r_early_rst),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_reset_req~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ociram_reset_req.extended_lut = "off";
defparam ociram_reset_req.lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam ociram_reset_req.shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[0]~0 (
	.dataa(!MonDReg_0),
	.datab(!\jtag_ram_access~q ),
	.datac(!writedata_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[0]~0 .extended_lut = "off";
defparam \ociram_wr_data[0]~0 .lut_mask = 64'h4747474747474747;
defparam \ociram_wr_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[0]~0 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[2]~q ),
	.datac(!address_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[0]~0 .extended_lut = "off";
defparam \ociram_addr[0]~0 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[1]~1 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(!address_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[1]~1 .extended_lut = "off";
defparam \ociram_addr[1]~1 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[2]~2 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[4]~q ),
	.datac(!address_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[2]~2 .extended_lut = "off";
defparam \ociram_addr[2]~2 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[3]~3 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[5]~q ),
	.datac(!address_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[3]~3 .extended_lut = "off";
defparam \ociram_addr[3]~3 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[4]~4 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[6]~q ),
	.datac(!address_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[4]~4 .extended_lut = "off";
defparam \ociram_addr[4]~4 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[5]~5 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[7]~q ),
	.datac(!address_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[5]~5 .extended_lut = "off";
defparam \ociram_addr[5]~5 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[6]~6 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[8]~q ),
	.datac(!address_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[6]~6 .extended_lut = "off";
defparam \ociram_addr[6]~6 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[7]~7 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[9]~q ),
	.datac(!address_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[7]~7 .extended_lut = "off";
defparam \ociram_addr[7]~7 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[0]~0 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[0]~0 .extended_lut = "off";
defparam \ociram_byteenable[0]~0 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[1]~1 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_1),
	.datac(!writedata_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[1]~1 .extended_lut = "off";
defparam \ociram_wr_data[1]~1 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \jtag_ram_wr~0 (
	.dataa(!take_action_ocimem_a),
	.datab(!jdo_35),
	.datac(!\Add0~1_sumout ),
	.datad(!\jtag_ram_wr~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_ram_wr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_ram_wr~0 .extended_lut = "off";
defparam \jtag_ram_wr~0 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \jtag_ram_wr~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[2]~2 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_2),
	.datac(!writedata_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[2]~2 .extended_lut = "off";
defparam \ociram_wr_data[2]~2 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[22]~3 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_22),
	.datac(!writedata_22),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[22]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[22]~3 .extended_lut = "off";
defparam \ociram_wr_data[22]~3 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[22]~3 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[2]~1 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[2]~1 .extended_lut = "off";
defparam \ociram_byteenable[2]~1 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[23]~4 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_23),
	.datac(!writedata_23),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[23]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[23]~4 .extended_lut = "off";
defparam \ociram_wr_data[23]~4 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[23]~4 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[24]~5 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_24),
	.datac(!writedata_24),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[24]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[24]~5 .extended_lut = "off";
defparam \ociram_wr_data[24]~5 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[24]~5 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[3]~2 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[3]~2 .extended_lut = "off";
defparam \ociram_byteenable[3]~2 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[25]~6 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_25),
	.datac(!writedata_25),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[25]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[25]~6 .extended_lut = "off";
defparam \ociram_wr_data[25]~6 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[25]~6 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[26]~7 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_26),
	.datac(!writedata_26),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[26]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[26]~7 .extended_lut = "off";
defparam \ociram_wr_data[26]~7 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[26]~7 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[11]~8 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_11),
	.datac(!writedata_11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[11]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[11]~8 .extended_lut = "off";
defparam \ociram_wr_data[11]~8 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[11]~8 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[1]~3 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[1]~3 .extended_lut = "off";
defparam \ociram_byteenable[1]~3 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[1]~3 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[12]~9 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_12),
	.datac(!writedata_12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[12]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[12]~9 .extended_lut = "off";
defparam \ociram_wr_data[12]~9 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[12]~9 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[13]~10 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_13),
	.datac(!writedata_13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[13]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[13]~10 .extended_lut = "off";
defparam \ociram_wr_data[13]~10 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[13]~10 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[14]~11 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_14),
	.datac(!writedata_14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[14]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[14]~11 .extended_lut = "off";
defparam \ociram_wr_data[14]~11 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[14]~11 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[15]~12 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_15),
	.datac(!writedata_15),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[15]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[15]~12 .extended_lut = "off";
defparam \ociram_wr_data[15]~12 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[15]~12 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[16]~13 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_16),
	.datac(!writedata_16),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[16]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[16]~13 .extended_lut = "off";
defparam \ociram_wr_data[16]~13 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[16]~13 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[3]~14 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_3),
	.datac(!writedata_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[3]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[3]~14 .extended_lut = "off";
defparam \ociram_wr_data[3]~14 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[3]~14 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[4]~15 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_4),
	.datac(!writedata_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[4]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[4]~15 .extended_lut = "off";
defparam \ociram_wr_data[4]~15 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[4]~15 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[5]~16 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_5),
	.datac(!writedata_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[5]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[5]~16 .extended_lut = "off";
defparam \ociram_wr_data[5]~16 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[5]~16 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[8]~17 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_8),
	.datac(!writedata_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[8]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[8]~17 .extended_lut = "off";
defparam \ociram_wr_data[8]~17 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[8]~17 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[10]~18 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_10),
	.datac(!writedata_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[10]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[10]~18 .extended_lut = "off";
defparam \ociram_wr_data[10]~18 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[10]~18 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[17]~19 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_17),
	.datac(!writedata_17),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[17]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[17]~19 .extended_lut = "off";
defparam \ociram_wr_data[17]~19 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[17]~19 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[9]~20 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_9),
	.datac(!writedata_9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[9]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[9]~20 .extended_lut = "off";
defparam \ociram_wr_data[9]~20 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[9]~20 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[18]~21 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_18),
	.datac(!writedata_18),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[18]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[18]~21 .extended_lut = "off";
defparam \ociram_wr_data[18]~21 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[18]~21 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[19]~22 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_19),
	.datac(!writedata_19),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[19]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[19]~22 .extended_lut = "off";
defparam \ociram_wr_data[19]~22 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[19]~22 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[20]~23 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_20),
	.datac(!writedata_20),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[20]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[20]~23 .extended_lut = "off";
defparam \ociram_wr_data[20]~23 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[20]~23 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[21]~24 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_21),
	.datac(!writedata_21),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[21]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[21]~24 .extended_lut = "off";
defparam \ociram_wr_data[21]~24 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[21]~24 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[6]~25 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_6),
	.datac(!writedata_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[6]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[6]~25 .extended_lut = "off";
defparam \ociram_wr_data[6]~25 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[6]~25 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[7]~26 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_7),
	.datac(!writedata_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[7]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[7]~26 .extended_lut = "off";
defparam \ociram_wr_data[7]~26 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[7]~26 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[27]~27 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_27),
	.datac(!writedata_27),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[27]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[27]~27 .extended_lut = "off";
defparam \ociram_wr_data[27]~27 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[27]~27 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[28]~28 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_28),
	.datac(!writedata_28),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[28]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[28]~28 .extended_lut = "off";
defparam \ociram_wr_data[28]~28 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[28]~28 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[29]~29 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_29),
	.datac(!writedata_29),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[29]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[29]~29 .extended_lut = "off";
defparam \ociram_wr_data[29]~29 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[29]~29 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[30]~30 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_30),
	.datac(!writedata_30),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[30]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[30]~30 .extended_lut = "off";
defparam \ociram_wr_data[30]~30 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[30]~30 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[31]~31 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_31),
	.datac(!writedata_31),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[31]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[31]~31 .extended_lut = "off";
defparam \ociram_wr_data[31]~31 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[31]~31 .shared_arith = "off";

dffeas \MonDReg[1] (
	.clk(clk_clk),
	.d(jdo_4),
	.asdata(q_a_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_1),
	.prn(vcc));
defparam \MonDReg[1] .is_wysiwyg = "true";
defparam \MonDReg[1] .power_up = "low";

dffeas \MonDReg[2] (
	.clk(clk_clk),
	.d(jdo_5),
	.asdata(q_a_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_2),
	.prn(vcc));
defparam \MonDReg[2] .is_wysiwyg = "true";
defparam \MonDReg[2] .power_up = "low";

dffeas \MonDReg[3] (
	.clk(clk_clk),
	.d(jdo_6),
	.asdata(q_a_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_3),
	.prn(vcc));
defparam \MonDReg[3] .is_wysiwyg = "true";
defparam \MonDReg[3] .power_up = "low";

dffeas \MonDReg[16] (
	.clk(clk_clk),
	.d(jdo_19),
	.asdata(q_a_16),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_16),
	.prn(vcc));
defparam \MonDReg[16] .is_wysiwyg = "true";
defparam \MonDReg[16] .power_up = "low";

dffeas \MonDReg[24] (
	.clk(clk_clk),
	.d(jdo_27),
	.asdata(q_a_24),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_24),
	.prn(vcc));
defparam \MonDReg[24] .is_wysiwyg = "true";
defparam \MonDReg[24] .power_up = "low";

dffeas \MonDReg[25] (
	.clk(clk_clk),
	.d(jdo_28),
	.asdata(q_a_25),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_25),
	.prn(vcc));
defparam \MonDReg[25] .is_wysiwyg = "true";
defparam \MonDReg[25] .power_up = "low";

dffeas \MonDReg[27] (
	.clk(clk_clk),
	.d(jdo_30),
	.asdata(q_a_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_27),
	.prn(vcc));
defparam \MonDReg[27] .is_wysiwyg = "true";
defparam \MonDReg[27] .power_up = "low";

dffeas \MonDReg[26] (
	.clk(clk_clk),
	.d(jdo_29),
	.asdata(q_a_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_26),
	.prn(vcc));
defparam \MonDReg[26] .is_wysiwyg = "true";
defparam \MonDReg[26] .power_up = "low";

dffeas \MonDReg[22] (
	.clk(clk_clk),
	.d(jdo_25),
	.asdata(q_a_22),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_22),
	.prn(vcc));
defparam \MonDReg[22] .is_wysiwyg = "true";
defparam \MonDReg[22] .power_up = "low";

dffeas \MonDReg[20] (
	.clk(clk_clk),
	.d(jdo_23),
	.asdata(q_a_20),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_20),
	.prn(vcc));
defparam \MonDReg[20] .is_wysiwyg = "true";
defparam \MonDReg[20] .power_up = "low";

dffeas \MonDReg[19] (
	.clk(clk_clk),
	.d(jdo_22),
	.asdata(q_a_19),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_19),
	.prn(vcc));
defparam \MonDReg[19] .is_wysiwyg = "true";
defparam \MonDReg[19] .power_up = "low";

dffeas \MonDReg[23] (
	.clk(clk_clk),
	.d(jdo_26),
	.asdata(q_a_23),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_23),
	.prn(vcc));
defparam \MonDReg[23] .is_wysiwyg = "true";
defparam \MonDReg[23] .power_up = "low";

dffeas \MonDReg[11] (
	.clk(clk_clk),
	.d(jdo_14),
	.asdata(q_a_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_11),
	.prn(vcc));
defparam \MonDReg[11] .is_wysiwyg = "true";
defparam \MonDReg[11] .power_up = "low";

dffeas \MonDReg[13] (
	.clk(clk_clk),
	.d(jdo_16),
	.asdata(q_a_13),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_13),
	.prn(vcc));
defparam \MonDReg[13] .is_wysiwyg = "true";
defparam \MonDReg[13] .power_up = "low";

dffeas \MonDReg[14] (
	.clk(clk_clk),
	.d(jdo_17),
	.asdata(q_a_14),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_14),
	.prn(vcc));
defparam \MonDReg[14] .is_wysiwyg = "true";
defparam \MonDReg[14] .power_up = "low";

dffeas \MonDReg[10] (
	.clk(clk_clk),
	.d(jdo_13),
	.asdata(q_a_10),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_10),
	.prn(vcc));
defparam \MonDReg[10] .is_wysiwyg = "true";
defparam \MonDReg[10] .power_up = "low";

dffeas \MonDReg[17] (
	.clk(clk_clk),
	.d(jdo_20),
	.asdata(q_a_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_17),
	.prn(vcc));
defparam \MonDReg[17] .is_wysiwyg = "true";
defparam \MonDReg[17] .power_up = "low";

dffeas \MonDReg[9] (
	.clk(clk_clk),
	.d(jdo_12),
	.asdata(q_a_9),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_9),
	.prn(vcc));
defparam \MonDReg[9] .is_wysiwyg = "true";
defparam \MonDReg[9] .power_up = "low";

dffeas \MonDReg[21] (
	.clk(clk_clk),
	.d(jdo_24),
	.asdata(q_a_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_21),
	.prn(vcc));
defparam \MonDReg[21] .is_wysiwyg = "true";
defparam \MonDReg[21] .power_up = "low";

dffeas \MonDReg[6] (
	.clk(clk_clk),
	.d(jdo_9),
	.asdata(q_a_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_6),
	.prn(vcc));
defparam \MonDReg[6] .is_wysiwyg = "true";
defparam \MonDReg[6] .power_up = "low";

dffeas \MonDReg[7] (
	.clk(clk_clk),
	.d(jdo_10),
	.asdata(q_a_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_7),
	.prn(vcc));
defparam \MonDReg[7] .is_wysiwyg = "true";
defparam \MonDReg[7] .power_up = "low";

dffeas \MonDReg[28] (
	.clk(clk_clk),
	.d(jdo_31),
	.asdata(q_a_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_28),
	.prn(vcc));
defparam \MonDReg[28] .is_wysiwyg = "true";
defparam \MonDReg[28] .power_up = "low";

dffeas \MonDReg[30] (
	.clk(clk_clk),
	.d(jdo_33),
	.asdata(q_a_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_30),
	.prn(vcc));
defparam \MonDReg[30] .is_wysiwyg = "true";
defparam \MonDReg[30] .power_up = "low";

dffeas \MonDReg[31] (
	.clk(clk_clk),
	.d(jdo_34),
	.asdata(q_a_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[11]~3_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_31),
	.prn(vcc));
defparam \MonDReg[31] .is_wysiwyg = "true";
defparam \MonDReg[31] .power_up = "low";

dffeas waitrequest(
	.clk(clk_clk),
	.d(\waitrequest~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest1),
	.prn(vcc));
defparam waitrequest.is_wysiwyg = "true";
defparam waitrequest.power_up = "low";

dffeas \MonDReg[0] (
	.clk(clk_clk),
	.d(\MonDReg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_0),
	.prn(vcc));
defparam \MonDReg[0] .is_wysiwyg = "true";
defparam \MonDReg[0] .power_up = "low";

dffeas \MonDReg[4] (
	.clk(clk_clk),
	.d(\MonDReg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_4),
	.prn(vcc));
defparam \MonDReg[4] .is_wysiwyg = "true";
defparam \MonDReg[4] .power_up = "low";

dffeas \MonDReg[12] (
	.clk(clk_clk),
	.d(\MonDReg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_12),
	.prn(vcc));
defparam \MonDReg[12] .is_wysiwyg = "true";
defparam \MonDReg[12] .power_up = "low";

dffeas \MonDReg[15] (
	.clk(clk_clk),
	.d(\MonDReg[15]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[15]~6_combout ),
	.q(MonDReg_15),
	.prn(vcc));
defparam \MonDReg[15] .is_wysiwyg = "true";
defparam \MonDReg[15] .power_up = "low";

dffeas \MonDReg[5] (
	.clk(clk_clk),
	.d(\MonDReg~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_5),
	.prn(vcc));
defparam \MonDReg[5] .is_wysiwyg = "true";
defparam \MonDReg[5] .power_up = "low";

dffeas \MonDReg[8] (
	.clk(clk_clk),
	.d(\MonDReg[8]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[15]~6_combout ),
	.q(MonDReg_8),
	.prn(vcc));
defparam \MonDReg[8] .is_wysiwyg = "true";
defparam \MonDReg[8] .power_up = "low";

dffeas \MonDReg[18] (
	.clk(clk_clk),
	.d(\MonDReg~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_18),
	.prn(vcc));
defparam \MonDReg[18] .is_wysiwyg = "true";
defparam \MonDReg[18] .power_up = "low";

dffeas \MonDReg[29] (
	.clk(clk_clk),
	.d(\MonDReg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_29),
	.prn(vcc));
defparam \MonDReg[29] .is_wysiwyg = "true";
defparam \MonDReg[29] .power_up = "low";

cyclonev_lcell_comb \Add0~1_wirecell (
	.dataa(!\Add0~1_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1_wirecell .extended_lut = "off";
defparam \Add0~1_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \Add0~1_wirecell .shared_arith = "off";

dffeas \MonAReg[10] (
	.clk(clk_clk),
	.d(\Add0~1_wirecell_combout ),
	.asdata(jdo_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[10]~q ),
	.prn(vcc));
defparam \MonAReg[10] .is_wysiwyg = "true";
defparam \MonAReg[10] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \MonAReg[2] (
	.clk(clk_clk),
	.d(\Add0~5_sumout ),
	.asdata(jdo_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[2]~q ),
	.prn(vcc));
defparam \MonAReg[2] .is_wysiwyg = "true";
defparam \MonAReg[2] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \MonAReg[3] (
	.clk(clk_clk),
	.d(\Add0~13_sumout ),
	.asdata(jdo_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[3]~q ),
	.prn(vcc));
defparam \MonAReg[3] .is_wysiwyg = "true";
defparam \MonAReg[3] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \MonAReg[4] (
	.clk(clk_clk),
	.d(\Add0~9_sumout ),
	.asdata(jdo_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[4]~q ),
	.prn(vcc));
defparam \MonAReg[4] .is_wysiwyg = "true";
defparam \MonAReg[4] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \MonAReg[5] (
	.clk(clk_clk),
	.d(\Add0~21_sumout ),
	.asdata(jdo_29),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[5]~q ),
	.prn(vcc));
defparam \MonAReg[5] .is_wysiwyg = "true";
defparam \MonAReg[5] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \MonAReg[6] (
	.clk(clk_clk),
	.d(\Add0~25_sumout ),
	.asdata(jdo_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[6]~q ),
	.prn(vcc));
defparam \MonAReg[6] .is_wysiwyg = "true";
defparam \MonAReg[6] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \MonAReg[7] (
	.clk(clk_clk),
	.d(\Add0~29_sumout ),
	.asdata(jdo_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[7]~q ),
	.prn(vcc));
defparam \MonAReg[7] .is_wysiwyg = "true";
defparam \MonAReg[7] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \MonAReg[8] (
	.clk(clk_clk),
	.d(\Add0~33_sumout ),
	.asdata(jdo_32),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[8]~q ),
	.prn(vcc));
defparam \MonAReg[8] .is_wysiwyg = "true";
defparam \MonAReg[8] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \MonAReg[9] (
	.clk(clk_clk),
	.d(\Add0~17_sumout ),
	.asdata(jdo_33),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[9]~q ),
	.prn(vcc));
defparam \MonAReg[9] .is_wysiwyg = "true";
defparam \MonAReg[9] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \jtag_ram_rd~0 (
	.dataa(!take_action_ocimem_a1),
	.datab(!jdo_34),
	.datac(!jdo_17),
	.datad(!\Add0~1_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_ram_rd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_ram_rd~0 .extended_lut = "off";
defparam \jtag_ram_rd~0 .lut_mask = 64'hD1FFD1FFD1FFD1FF;
defparam \jtag_ram_rd~0 .shared_arith = "off";

dffeas jtag_ram_rd(
	.clk(clk_clk),
	.d(\jtag_ram_rd~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!take_action_ocimem_b),
	.q(\jtag_ram_rd~q ),
	.prn(vcc));
defparam jtag_ram_rd.is_wysiwyg = "true";
defparam jtag_ram_rd.power_up = "low";

dffeas jtag_ram_rd_d1(
	.clk(clk_clk),
	.d(\jtag_ram_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_rd_d1~q ),
	.prn(vcc));
defparam jtag_ram_rd_d1.is_wysiwyg = "true";
defparam jtag_ram_rd_d1.power_up = "low";

cyclonev_lcell_comb \MonDReg[11]~3 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[11]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[11]~3 .extended_lut = "off";
defparam \MonDReg[11]~3 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \MonDReg[11]~3 .shared_arith = "off";

dffeas jtag_rd(
	.clk(clk_clk),
	.d(take_action_ocimem_a1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!take_action_ocimem_b),
	.q(\jtag_rd~q ),
	.prn(vcc));
defparam jtag_rd.is_wysiwyg = "true";
defparam jtag_rd.power_up = "low";

dffeas jtag_rd_d1(
	.clk(clk_clk),
	.d(\jtag_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_rd_d1~q ),
	.prn(vcc));
defparam jtag_rd_d1.is_wysiwyg = "true";
defparam jtag_rd_d1.power_up = "low";

cyclonev_lcell_comb \MonDReg[0]~2 (
	.dataa(!ir_1),
	.datab(!ir_0),
	.datac(!enable_action_strobe),
	.datad(!jdo_35),
	.datae(!\jtag_rd_d1~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[0]~2 .extended_lut = "off";
defparam \MonDReg[0]~2 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \MonDReg[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \jtag_ram_access~0 (
	.dataa(!take_action_ocimem_a),
	.datab(!jdo_35),
	.datac(!jdo_34),
	.datad(!jdo_17),
	.datae(!\Add0~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_ram_access~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_ram_access~0 .extended_lut = "off";
defparam \jtag_ram_access~0 .lut_mask = 64'hFF7DFFFFFF7DFFFF;
defparam \jtag_ram_access~0 .shared_arith = "off";

dffeas jtag_ram_access(
	.clk(clk_clk),
	.d(\jtag_ram_access~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_access~q ),
	.prn(vcc));
defparam jtag_ram_access.is_wysiwyg = "true";
defparam jtag_ram_access.power_up = "low";

cyclonev_lcell_comb \waitrequest~0 (
	.dataa(!address_8),
	.datab(!\jtag_ram_access~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\waitrequest~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \waitrequest~0 .extended_lut = "off";
defparam \waitrequest~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \waitrequest~0 .shared_arith = "off";

cyclonev_lcell_comb \avalon_ociram_readdata_ready~0 (
	.dataa(!waitrequest1),
	.datab(!write),
	.datac(!\waitrequest~0_combout ),
	.datad(!read),
	.datae(!\avalon_ociram_readdata_ready~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\avalon_ociram_readdata_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \avalon_ociram_readdata_ready~0 .extended_lut = "off";
defparam \avalon_ociram_readdata_ready~0 .lut_mask = 64'hD1FFFFFFD1FFFFFF;
defparam \avalon_ociram_readdata_ready~0 .shared_arith = "off";

dffeas avalon_ociram_readdata_ready(
	.clk(clk_clk),
	.d(\avalon_ociram_readdata_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\avalon_ociram_readdata_ready~q ),
	.prn(vcc));
defparam avalon_ociram_readdata_ready.is_wysiwyg = "true";
defparam avalon_ociram_readdata_ready.power_up = "low";

cyclonev_lcell_comb \waitrequest~1 (
	.dataa(!waitrequest1),
	.datab(!write),
	.datac(!\waitrequest~0_combout ),
	.datad(!read),
	.datae(!\avalon_ociram_readdata_ready~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\waitrequest~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \waitrequest~1 .extended_lut = "off";
defparam \waitrequest~1 .lut_mask = 64'hFFFFBF8FFFFFBF8F;
defparam \waitrequest~1 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~0 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonAReg[2]~q ),
	.datac(!\MonAReg[4]~q ),
	.datad(!\MonAReg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~0 .extended_lut = "off";
defparam \MonDReg~0 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \MonDReg~0 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~1 (
	.dataa(!take_action_ocimem_b),
	.datab(!jdo_3),
	.datac(!\jtag_ram_rd_d1~q ),
	.datad(!q_a_0),
	.datae(!\MonDReg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~1 .extended_lut = "off";
defparam \MonDReg~1 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~1 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~4 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonDReg~0_combout ),
	.datad(!q_a_4),
	.datae(!jdo_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~4 .extended_lut = "off";
defparam \MonDReg~4 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~4 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~5 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonDReg~0_combout ),
	.datad(!q_a_12),
	.datae(!jdo_15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~5 .extended_lut = "off";
defparam \MonDReg~5 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \MonDReg~5 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg[15]~20 (
	.dataa(!\MonAReg[4]~q ),
	.datab(!\MonAReg[2]~q ),
	.datac(!q_a_15),
	.datad(!jdo_18),
	.datae(!\jtag_ram_rd_d1~q ),
	.dataf(!take_action_ocimem_b),
	.datag(!\MonAReg[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[15]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[15]~20 .extended_lut = "on";
defparam \MonDReg[15]~20 .lut_mask = 64'hFF6FFFF6FF6FFFF6;
defparam \MonDReg[15]~20 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg[15]~6 (
	.dataa(!ir_1),
	.datab(!ir_0),
	.datac(!enable_action_strobe),
	.datad(!jdo_35),
	.datae(!\jtag_rd_d1~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[15]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[15]~6 .extended_lut = "off";
defparam \MonDReg[15]~6 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \MonDReg[15]~6 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~16 (
	.dataa(!\MonAReg[3]~q ),
	.datab(!\MonAReg[4]~q ),
	.datac(!q_a_5),
	.datad(!jdo_8),
	.datae(!\jtag_ram_rd_d1~q ),
	.dataf(!take_action_ocimem_b),
	.datag(!\MonAReg[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~16 .extended_lut = "on";
defparam \MonDReg~16 .lut_mask = 64'hFF7FFFF7FF7FFFF7;
defparam \MonDReg~16 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg[8]~7 (
	.dataa(!take_action_ocimem_b),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonAReg[2]~q ),
	.datad(!\MonAReg[4]~q ),
	.datae(!q_a_8),
	.dataf(!jdo_11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[8]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[8]~7 .extended_lut = "off";
defparam \MonDReg[8]~7 .lut_mask = 64'hFF6FFFFFFFFFFFFF;
defparam \MonDReg[8]~7 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~12 (
	.dataa(!\MonAReg[3]~q ),
	.datab(!\MonAReg[4]~q ),
	.datac(!q_a_18),
	.datad(!jdo_21),
	.datae(!\jtag_ram_rd_d1~q ),
	.dataf(!take_action_ocimem_b),
	.datag(!\MonAReg[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~12 .extended_lut = "on";
defparam \MonDReg~12 .lut_mask = 64'hFFBFFFFBFFBFFFFB;
defparam \MonDReg~12 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~8 (
	.dataa(!\MonAReg[3]~q ),
	.datab(!\MonAReg[4]~q ),
	.datac(!q_a_29),
	.datad(!jdo_32),
	.datae(!\jtag_ram_rd_d1~q ),
	.dataf(!take_action_ocimem_b),
	.datag(!\MonAReg[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~8 .extended_lut = "on";
defparam \MonDReg~8 .lut_mask = 64'hFFDFFFFDFFDFFFFD;
defparam \MonDReg~8 .shared_arith = "off";

endmodule

module niosLab2_niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_11,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_15,
	q_a_16,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_8,
	q_a_10,
	q_a_17,
	q_a_9,
	q_a_18,
	q_a_19,
	q_a_20,
	q_a_21,
	q_a_6,
	q_a_7,
	q_a_27,
	q_a_28,
	q_a_29,
	q_a_30,
	q_a_31,
	ociram_wr_en,
	ociram_reset_req,
	ociram_wr_data_0,
	ociram_addr_0,
	ociram_addr_1,
	ociram_addr_2,
	ociram_addr_3,
	ociram_addr_4,
	ociram_addr_5,
	ociram_addr_6,
	ociram_addr_7,
	ociram_byteenable_0,
	ociram_wr_data_1,
	ociram_wr_data_2,
	ociram_wr_data_22,
	ociram_byteenable_2,
	ociram_wr_data_23,
	ociram_wr_data_24,
	ociram_byteenable_3,
	ociram_wr_data_25,
	ociram_wr_data_26,
	ociram_wr_data_11,
	ociram_byteenable_1,
	ociram_wr_data_12,
	ociram_wr_data_13,
	ociram_wr_data_14,
	ociram_wr_data_15,
	ociram_wr_data_16,
	ociram_wr_data_3,
	ociram_wr_data_4,
	ociram_wr_data_5,
	ociram_wr_data_8,
	ociram_wr_data_10,
	ociram_wr_data_17,
	ociram_wr_data_9,
	ociram_wr_data_18,
	ociram_wr_data_19,
	ociram_wr_data_20,
	ociram_wr_data_21,
	ociram_wr_data_6,
	ociram_wr_data_7,
	ociram_wr_data_27,
	ociram_wr_data_28,
	ociram_wr_data_29,
	ociram_wr_data_30,
	ociram_wr_data_31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_22;
output 	q_a_23;
output 	q_a_24;
output 	q_a_25;
output 	q_a_26;
output 	q_a_11;
output 	q_a_12;
output 	q_a_13;
output 	q_a_14;
output 	q_a_15;
output 	q_a_16;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_8;
output 	q_a_10;
output 	q_a_17;
output 	q_a_9;
output 	q_a_18;
output 	q_a_19;
output 	q_a_20;
output 	q_a_21;
output 	q_a_6;
output 	q_a_7;
output 	q_a_27;
output 	q_a_28;
output 	q_a_29;
output 	q_a_30;
output 	q_a_31;
input 	ociram_wr_en;
input 	ociram_reset_req;
input 	ociram_wr_data_0;
input 	ociram_addr_0;
input 	ociram_addr_1;
input 	ociram_addr_2;
input 	ociram_addr_3;
input 	ociram_addr_4;
input 	ociram_addr_5;
input 	ociram_addr_6;
input 	ociram_addr_7;
input 	ociram_byteenable_0;
input 	ociram_wr_data_1;
input 	ociram_wr_data_2;
input 	ociram_wr_data_22;
input 	ociram_byteenable_2;
input 	ociram_wr_data_23;
input 	ociram_wr_data_24;
input 	ociram_byteenable_3;
input 	ociram_wr_data_25;
input 	ociram_wr_data_26;
input 	ociram_wr_data_11;
input 	ociram_byteenable_1;
input 	ociram_wr_data_12;
input 	ociram_wr_data_13;
input 	ociram_wr_data_14;
input 	ociram_wr_data_15;
input 	ociram_wr_data_16;
input 	ociram_wr_data_3;
input 	ociram_wr_data_4;
input 	ociram_wr_data_5;
input 	ociram_wr_data_8;
input 	ociram_wr_data_10;
input 	ociram_wr_data_17;
input 	ociram_wr_data_9;
input 	ociram_wr_data_18;
input 	ociram_wr_data_19;
input 	ociram_wr_data_20;
input 	ociram_wr_data_21;
input 	ociram_wr_data_6;
input 	ociram_wr_data_7;
input 	ociram_wr_data_27;
input 	ociram_wr_data_28;
input 	ociram_wr_data_29;
input 	ociram_wr_data_30;
input 	ociram_wr_data_31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosLab2_altsyncram_1 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.wren_a(ociram_wr_en),
	.clocken0(ociram_reset_req),
	.data_a({ociram_wr_data_31,ociram_wr_data_30,ociram_wr_data_29,ociram_wr_data_28,ociram_wr_data_27,ociram_wr_data_26,ociram_wr_data_25,ociram_wr_data_24,ociram_wr_data_23,ociram_wr_data_22,ociram_wr_data_21,ociram_wr_data_20,ociram_wr_data_19,ociram_wr_data_18,ociram_wr_data_17,
ociram_wr_data_16,ociram_wr_data_15,ociram_wr_data_14,ociram_wr_data_13,ociram_wr_data_12,ociram_wr_data_11,ociram_wr_data_10,ociram_wr_data_9,ociram_wr_data_8,ociram_wr_data_7,ociram_wr_data_6,ociram_wr_data_5,ociram_wr_data_4,ociram_wr_data_3,ociram_wr_data_2,
ociram_wr_data_1,ociram_wr_data_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,ociram_addr_7,ociram_addr_6,ociram_addr_5,ociram_addr_4,ociram_addr_3,ociram_addr_2,ociram_addr_1,ociram_addr_0}),
	.byteena_a({ociram_byteenable_3,ociram_byteenable_2,ociram_byteenable_1,ociram_byteenable_0}),
	.clock0(clk_clk));

endmodule

module niosLab2_altsyncram_1 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosLab2_altsyncram_qid1 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module niosLab2_altsyncram_qid1 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 8;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 255;
defparam ram_block1a22.port_a_logical_ram_depth = 256;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 8;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 255;
defparam ram_block1a23.port_a_logical_ram_depth = 256;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 8;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 255;
defparam ram_block1a24.port_a_logical_ram_depth = 256;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 8;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 255;
defparam ram_block1a25.port_a_logical_ram_depth = 256;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 8;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 255;
defparam ram_block1a26.port_a_logical_ram_depth = 256;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 8;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 255;
defparam ram_block1a20.port_a_logical_ram_depth = 256;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 8;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 255;
defparam ram_block1a21.port_a_logical_ram_depth = 256;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 8;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 255;
defparam ram_block1a27.port_a_logical_ram_depth = 256;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 8;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 255;
defparam ram_block1a28.port_a_logical_ram_depth = 256;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 8;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 255;
defparam ram_block1a29.port_a_logical_ram_depth = 256;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a29.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 8;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 255;
defparam ram_block1a30.port_a_logical_ram_depth = 256;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_nios2_oci:the_niosLab2_nios2_gen2_0_cpu_nios2_oci|niosLab2_nios2_gen2_0_cpu_nios2_ocimem:the_niosLab2_nios2_gen2_0_cpu_nios2_ocimem|niosLab2_nios2_gen2_0_cpu_ociram_sp_ram_module:niosLab2_nios2_gen2_0_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_qid1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 8;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 255;
defparam ram_block1a31.port_a_logical_ram_depth = 256;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a31.ram_block_type = "auto";

endmodule

module niosLab2_niosLab2_nios2_gen2_0_cpu_register_bank_a_module (
	q_b_4,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_3,
	q_b_2,
	D_iw_27,
	D_iw_28,
	D_iw_29,
	D_iw_30,
	D_iw_31,
	q_b_25,
	q_b_27,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_18,
	q_b_17,
	q_b_1,
	q_b_26,
	q_b_31,
	q_b_30,
	q_b_0,
	q_b_28,
	q_b_29,
	W_rf_wr_data_0,
	W_rf_wren,
	R_dst_regnum_0,
	R_dst_regnum_1,
	R_dst_regnum_2,
	R_dst_regnum_3,
	R_dst_regnum_4,
	W_rf_wr_data_1,
	W_rf_wr_data_2,
	W_rf_wr_data_3,
	W_rf_wr_data_4,
	W_rf_wr_data_5,
	W_rf_wr_data_11,
	W_rf_wr_data_10,
	W_rf_wr_data_9,
	W_rf_wr_data_8,
	W_rf_wr_data_7,
	W_rf_wr_data_6,
	W_rf_wr_data_12,
	W_rf_wr_data_13,
	W_rf_wr_data_14,
	W_rf_wr_data_15,
	W_rf_wr_data_16,
	W_rf_wr_data_25,
	W_rf_wr_data_27,
	W_rf_wr_data_19,
	W_rf_wr_data_20,
	W_rf_wr_data_21,
	W_rf_wr_data_22,
	W_rf_wr_data_23,
	W_rf_wr_data_24,
	W_rf_wr_data_18,
	W_rf_wr_data_17,
	W_rf_wr_data_26,
	W_rf_wr_data_31,
	W_rf_wr_data_30,
	W_rf_wr_data_28,
	W_rf_wr_data_29,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_4;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_3;
output 	q_b_2;
input 	D_iw_27;
input 	D_iw_28;
input 	D_iw_29;
input 	D_iw_30;
input 	D_iw_31;
output 	q_b_25;
output 	q_b_27;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_24;
output 	q_b_18;
output 	q_b_17;
output 	q_b_1;
output 	q_b_26;
output 	q_b_31;
output 	q_b_30;
output 	q_b_0;
output 	q_b_28;
output 	q_b_29;
input 	W_rf_wr_data_0;
input 	W_rf_wren;
input 	R_dst_regnum_0;
input 	R_dst_regnum_1;
input 	R_dst_regnum_2;
input 	R_dst_regnum_3;
input 	R_dst_regnum_4;
input 	W_rf_wr_data_1;
input 	W_rf_wr_data_2;
input 	W_rf_wr_data_3;
input 	W_rf_wr_data_4;
input 	W_rf_wr_data_5;
input 	W_rf_wr_data_11;
input 	W_rf_wr_data_10;
input 	W_rf_wr_data_9;
input 	W_rf_wr_data_8;
input 	W_rf_wr_data_7;
input 	W_rf_wr_data_6;
input 	W_rf_wr_data_12;
input 	W_rf_wr_data_13;
input 	W_rf_wr_data_14;
input 	W_rf_wr_data_15;
input 	W_rf_wr_data_16;
input 	W_rf_wr_data_25;
input 	W_rf_wr_data_27;
input 	W_rf_wr_data_19;
input 	W_rf_wr_data_20;
input 	W_rf_wr_data_21;
input 	W_rf_wr_data_22;
input 	W_rf_wr_data_23;
input 	W_rf_wr_data_24;
input 	W_rf_wr_data_18;
input 	W_rf_wr_data_17;
input 	W_rf_wr_data_26;
input 	W_rf_wr_data_31;
input 	W_rf_wr_data_30;
input 	W_rf_wr_data_28;
input 	W_rf_wr_data_29;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosLab2_altsyncram_2 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_b({D_iw_31,D_iw_30,D_iw_29,D_iw_28,D_iw_27}),
	.data_a({W_rf_wr_data_31,W_rf_wr_data_30,W_rf_wr_data_29,W_rf_wr_data_28,W_rf_wr_data_27,W_rf_wr_data_26,W_rf_wr_data_25,W_rf_wr_data_24,W_rf_wr_data_23,W_rf_wr_data_22,W_rf_wr_data_21,W_rf_wr_data_20,W_rf_wr_data_19,W_rf_wr_data_18,W_rf_wr_data_17,W_rf_wr_data_16,W_rf_wr_data_15,
W_rf_wr_data_14,W_rf_wr_data_13,W_rf_wr_data_12,W_rf_wr_data_11,W_rf_wr_data_10,W_rf_wr_data_9,W_rf_wr_data_8,W_rf_wr_data_7,W_rf_wr_data_6,W_rf_wr_data_5,W_rf_wr_data_4,W_rf_wr_data_3,W_rf_wr_data_2,W_rf_wr_data_1,W_rf_wr_data_0}),
	.wren_a(W_rf_wren),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,R_dst_regnum_4,R_dst_regnum_3,R_dst_regnum_2,R_dst_regnum_1,R_dst_regnum_0}),
	.clock0(clk_clk));

endmodule

module niosLab2_altsyncram_2 (
	q_b,
	address_b,
	data_a,
	wren_a,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[4:0] address_b;
input 	[31:0] data_a;
input 	wren_a;
input 	[12:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosLab2_altsyncram_msi1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.wren_a(wren_a),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module niosLab2_altsyncram_msi1 (
	q_b,
	address_b,
	data_a,
	wren_a,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[4:0] address_b;
input 	[31:0] data_a;
input 	wren_a;
input 	[4:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_a_module:niosLab2_nios2_gen2_0_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

endmodule

module niosLab2_niosLab2_nios2_gen2_0_cpu_register_bank_b_module (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	D_iw_22,
	D_iw_23,
	D_iw_24,
	D_iw_25,
	D_iw_26,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_7,
	q_b_6,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_25,
	q_b_27,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_18,
	q_b_17,
	q_b_26,
	q_b_31,
	q_b_30,
	q_b_28,
	q_b_29,
	W_rf_wr_data_0,
	W_rf_wren,
	R_dst_regnum_0,
	R_dst_regnum_1,
	R_dst_regnum_2,
	R_dst_regnum_3,
	R_dst_regnum_4,
	W_rf_wr_data_1,
	W_rf_wr_data_2,
	W_rf_wr_data_3,
	W_rf_wr_data_4,
	W_rf_wr_data_5,
	W_rf_wr_data_11,
	W_rf_wr_data_10,
	W_rf_wr_data_9,
	W_rf_wr_data_8,
	W_rf_wr_data_7,
	W_rf_wr_data_6,
	W_rf_wr_data_12,
	W_rf_wr_data_13,
	W_rf_wr_data_14,
	W_rf_wr_data_15,
	W_rf_wr_data_16,
	W_rf_wr_data_25,
	W_rf_wr_data_27,
	W_rf_wr_data_19,
	W_rf_wr_data_20,
	W_rf_wr_data_21,
	W_rf_wr_data_22,
	W_rf_wr_data_23,
	W_rf_wr_data_24,
	W_rf_wr_data_18,
	W_rf_wr_data_17,
	W_rf_wr_data_26,
	W_rf_wr_data_31,
	W_rf_wr_data_30,
	W_rf_wr_data_28,
	W_rf_wr_data_29,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
input 	D_iw_22;
input 	D_iw_23;
input 	D_iw_24;
input 	D_iw_25;
input 	D_iw_26;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_7;
output 	q_b_6;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_25;
output 	q_b_27;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_24;
output 	q_b_18;
output 	q_b_17;
output 	q_b_26;
output 	q_b_31;
output 	q_b_30;
output 	q_b_28;
output 	q_b_29;
input 	W_rf_wr_data_0;
input 	W_rf_wren;
input 	R_dst_regnum_0;
input 	R_dst_regnum_1;
input 	R_dst_regnum_2;
input 	R_dst_regnum_3;
input 	R_dst_regnum_4;
input 	W_rf_wr_data_1;
input 	W_rf_wr_data_2;
input 	W_rf_wr_data_3;
input 	W_rf_wr_data_4;
input 	W_rf_wr_data_5;
input 	W_rf_wr_data_11;
input 	W_rf_wr_data_10;
input 	W_rf_wr_data_9;
input 	W_rf_wr_data_8;
input 	W_rf_wr_data_7;
input 	W_rf_wr_data_6;
input 	W_rf_wr_data_12;
input 	W_rf_wr_data_13;
input 	W_rf_wr_data_14;
input 	W_rf_wr_data_15;
input 	W_rf_wr_data_16;
input 	W_rf_wr_data_25;
input 	W_rf_wr_data_27;
input 	W_rf_wr_data_19;
input 	W_rf_wr_data_20;
input 	W_rf_wr_data_21;
input 	W_rf_wr_data_22;
input 	W_rf_wr_data_23;
input 	W_rf_wr_data_24;
input 	W_rf_wr_data_18;
input 	W_rf_wr_data_17;
input 	W_rf_wr_data_26;
input 	W_rf_wr_data_31;
input 	W_rf_wr_data_30;
input 	W_rf_wr_data_28;
input 	W_rf_wr_data_29;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosLab2_altsyncram_3 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_b({D_iw_26,D_iw_25,D_iw_24,D_iw_23,D_iw_22}),
	.data_a({W_rf_wr_data_31,W_rf_wr_data_30,W_rf_wr_data_29,W_rf_wr_data_28,W_rf_wr_data_27,W_rf_wr_data_26,W_rf_wr_data_25,W_rf_wr_data_24,W_rf_wr_data_23,W_rf_wr_data_22,W_rf_wr_data_21,W_rf_wr_data_20,W_rf_wr_data_19,W_rf_wr_data_18,W_rf_wr_data_17,W_rf_wr_data_16,W_rf_wr_data_15,
W_rf_wr_data_14,W_rf_wr_data_13,W_rf_wr_data_12,W_rf_wr_data_11,W_rf_wr_data_10,W_rf_wr_data_9,W_rf_wr_data_8,W_rf_wr_data_7,W_rf_wr_data_6,W_rf_wr_data_5,W_rf_wr_data_4,W_rf_wr_data_3,W_rf_wr_data_2,W_rf_wr_data_1,W_rf_wr_data_0}),
	.wren_a(W_rf_wren),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,R_dst_regnum_4,R_dst_regnum_3,R_dst_regnum_2,R_dst_regnum_1,R_dst_regnum_0}),
	.clock0(clk_clk));

endmodule

module niosLab2_altsyncram_3 (
	q_b,
	address_b,
	data_a,
	wren_a,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[4:0] address_b;
input 	[31:0] data_a;
input 	wren_a;
input 	[12:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosLab2_altsyncram_msi1_1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.wren_a(wren_a),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module niosLab2_altsyncram_msi1_1 (
	q_b,
	address_b,
	data_a,
	wren_a,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[4:0] address_b;
input 	[31:0] data_a;
input 	wren_a;
input 	[4:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "niosLab2_nios2_gen2_0:nios2_gen2_0|niosLab2_nios2_gen2_0_cpu:cpu|niosLab2_nios2_gen2_0_cpu_register_bank_b_module:niosLab2_nios2_gen2_0_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_msi1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

endmodule

module niosLab2_niosLab2_onchip_memory2_0 (
	q_a_0,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_11,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_15,
	q_a_16,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_8,
	q_a_10,
	q_a_17,
	q_a_9,
	q_a_18,
	q_a_19,
	q_a_20,
	q_a_21,
	q_a_6,
	q_a_7,
	q_a_27,
	q_a_28,
	q_a_29,
	q_a_30,
	q_a_31,
	always2,
	saved_grant_0,
	mem_used_1,
	src2_valid,
	src_valid,
	r_early_rst,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	src_data_32,
	src_payload1,
	src_data_34,
	src_payload2,
	src_payload3,
	src_data_35,
	src_payload4,
	src_payload5,
	src_payload6,
	src_data_33,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_22;
output 	q_a_23;
output 	q_a_24;
output 	q_a_25;
output 	q_a_26;
output 	q_a_11;
output 	q_a_12;
output 	q_a_13;
output 	q_a_14;
output 	q_a_15;
output 	q_a_16;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_8;
output 	q_a_10;
output 	q_a_17;
output 	q_a_9;
output 	q_a_18;
output 	q_a_19;
output 	q_a_20;
output 	q_a_21;
output 	q_a_6;
output 	q_a_7;
output 	q_a_27;
output 	q_a_28;
output 	q_a_29;
output 	q_a_30;
output 	q_a_31;
input 	always2;
input 	saved_grant_0;
input 	mem_used_1;
input 	src2_valid;
input 	src_valid;
input 	r_early_rst;
input 	src_payload;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_46;
input 	src_data_47;
input 	src_data_48;
input 	src_data_49;
input 	src_data_50;
input 	src_data_32;
input 	src_payload1;
input 	src_data_34;
input 	src_payload2;
input 	src_payload3;
input 	src_data_35;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_data_33;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wren~0_combout ;


niosLab2_altsyncram_4 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(r_early_rst),
	.wren_a(\wren~0_combout ),
	.data_a({src_payload31,src_payload30,src_payload29,src_payload28,src_payload27,src_payload5,src_payload4,src_payload3,src_payload2,src_payload1,src_payload24,src_payload23,src_payload22,src_payload21,src_payload19,src_payload11,src_payload10,src_payload9,src_payload8,src_payload7,
src_payload6,src_payload18,src_payload20,src_payload17,src_payload26,src_payload25,src_payload16,src_payload15,src_payload14,src_payload13,src_payload12,src_payload}),
	.address_a({src_data_50,src_data_49,src_data_48,src_data_47,src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.byteena_a({src_data_35,src_data_34,src_data_33,src_data_32}),
	.clock0(clk_clk));

cyclonev_lcell_comb \wren~0 (
	.dataa(!always2),
	.datab(!saved_grant_0),
	.datac(!mem_used_1),
	.datad(!src2_valid),
	.datae(!src_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wren~0 .extended_lut = "off";
defparam \wren~0 .lut_mask = 64'hFFFFFFEFFFFFFFEF;
defparam \wren~0 .shared_arith = "off";

endmodule

module niosLab2_altsyncram_4 (
	q_a,
	clocken0,
	wren_a,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	clocken0;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



niosLab2_altsyncram_ddn1 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module niosLab2_altsyncram_ddn1 (
	q_a,
	clocken0,
	wren_a,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	clocken0;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 13;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 8191;
defparam ram_block1a0.port_a_logical_ram_depth = 8192;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a0.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a0.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a0.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a22(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 13;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 8191;
defparam ram_block1a22.port_a_logical_ram_depth = 8192;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a22.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a22.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a22.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a23(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 13;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 8191;
defparam ram_block1a23.port_a_logical_ram_depth = 8192;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a24(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 13;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 8191;
defparam ram_block1a24.port_a_logical_ram_depth = 8192;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a24.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a24.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a24.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a25(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 13;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 8191;
defparam ram_block1a25.port_a_logical_ram_depth = 8192;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a25.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a25.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a25.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a26(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 13;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 8191;
defparam ram_block1a26.port_a_logical_ram_depth = 8192;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a26.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a26.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a26.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a11(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 13;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 8191;
defparam ram_block1a11.port_a_logical_ram_depth = 8192;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a11.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a11.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a11.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a12(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 13;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 8191;
defparam ram_block1a12.port_a_logical_ram_depth = 8192;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a12.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a12.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a12.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a13(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 13;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 8191;
defparam ram_block1a13.port_a_logical_ram_depth = 8192;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a13.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a13.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a13.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a14(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 13;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 8191;
defparam ram_block1a14.port_a_logical_ram_depth = 8192;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a14.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a14.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a14.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a15(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 13;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 8191;
defparam ram_block1a15.port_a_logical_ram_depth = 8192;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a16(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 13;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 8191;
defparam ram_block1a16.port_a_logical_ram_depth = 8192;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a16.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a16.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a16.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a1(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 13;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 8191;
defparam ram_block1a1.port_a_logical_ram_depth = 8192;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a1.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a1.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a1.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a2(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 13;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 8191;
defparam ram_block1a2.port_a_logical_ram_depth = 8192;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a2.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a2.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a2.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a3(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 13;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 8191;
defparam ram_block1a3.port_a_logical_ram_depth = 8192;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a3.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a3.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a3.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a4(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 13;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 8191;
defparam ram_block1a4.port_a_logical_ram_depth = 8192;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a4.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a4.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a4.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a5(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 13;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 8191;
defparam ram_block1a5.port_a_logical_ram_depth = 8192;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a5.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a5.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a5.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a8(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 13;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 8191;
defparam ram_block1a8.port_a_logical_ram_depth = 8192;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a8.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a8.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a8.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a10(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 13;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 8191;
defparam ram_block1a10.port_a_logical_ram_depth = 8192;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a17(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 13;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 8191;
defparam ram_block1a17.port_a_logical_ram_depth = 8192;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a17.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a17.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a17.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a9(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 13;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 8191;
defparam ram_block1a9.port_a_logical_ram_depth = 8192;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a9.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a9.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a9.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a18(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 13;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 8191;
defparam ram_block1a18.port_a_logical_ram_depth = 8192;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a18.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a18.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a18.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a19(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 13;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 8191;
defparam ram_block1a19.port_a_logical_ram_depth = 8192;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a19.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a19.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a19.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a20(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 13;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 8191;
defparam ram_block1a20.port_a_logical_ram_depth = 8192;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a20.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a20.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a20.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a21(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 13;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 8191;
defparam ram_block1a21.port_a_logical_ram_depth = 8192;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a21.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a21.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a21.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a6(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 13;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 8191;
defparam ram_block1a6.port_a_logical_ram_depth = 8192;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a6.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a6.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a6.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a7(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 13;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 8191;
defparam ram_block1a7.port_a_logical_ram_depth = 8192;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a7.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a7.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a7.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a27(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 13;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 8191;
defparam ram_block1a27.port_a_logical_ram_depth = 8192;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a27.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a27.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a27.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a28(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 13;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 8191;
defparam ram_block1a28.port_a_logical_ram_depth = 8192;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a28.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a28.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a28.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a29(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 13;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 8191;
defparam ram_block1a29.port_a_logical_ram_depth = 8192;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a29.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a29.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a29.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a30(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 13;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 8191;
defparam ram_block1a30.port_a_logical_ram_depth = 8192;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a30.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a30.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a30.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a31(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "niosLab2_onchip_memory2_0.hex";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "niosLab2_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_ddn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 13;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 8191;
defparam ram_block1a31.port_a_logical_ram_depth = 8192;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

endmodule

module niosLab2_niosLab2_pio_0 (
	W_alu_result_4,
	W_alu_result_3,
	W_alu_result_2,
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	writedata,
	reset_n,
	mem_used_1,
	Equal2,
	Equal21,
	rst1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	d_write,
	write_accepted,
	always0,
	always01,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_3;
input 	W_alu_result_2;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
input 	[31:0] writedata;
input 	reset_n;
input 	mem_used_1;
input 	Equal2;
input 	Equal21;
input 	rst1;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	d_write;
input 	write_accepted;
output 	always0;
output 	always01;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \always0~1_combout ;
wire \always0~2_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

cyclonev_lcell_comb \always0~3 (
	.dataa(!rst1),
	.datab(!wait_latency_counter_1),
	.datac(!W_alu_result_4),
	.datad(!Equal2),
	.datae(!Equal21),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always0),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~3 .extended_lut = "off";
defparam \always0~3 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \always0~3 .shared_arith = "off";

cyclonev_lcell_comb \always0~4 (
	.dataa(!mem_used_1),
	.datab(!rst1),
	.datac(!wait_latency_counter_1),
	.datad(!W_alu_result_4),
	.datae(!Equal2),
	.dataf(!Equal21),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always01),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~4 .extended_lut = "off";
defparam \always0~4 .lut_mask = 64'hFFFBFFFFFFFFFFFF;
defparam \always0~4 .shared_arith = "off";

cyclonev_lcell_comb \readdata[0]~0 (
	.dataa(!data_out_0),
	.datab(!W_alu_result_3),
	.datac(!W_alu_result_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0]~0 .extended_lut = "off";
defparam \readdata[0]~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \readdata[1]~1 (
	.dataa(!data_out_1),
	.datab(!W_alu_result_3),
	.datac(!W_alu_result_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[1]~1 .extended_lut = "off";
defparam \readdata[1]~1 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \readdata[2]~2 (
	.dataa(!data_out_2),
	.datab(!W_alu_result_3),
	.datac(!W_alu_result_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[2]~2 .extended_lut = "off";
defparam \readdata[2]~2 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \readdata[3]~3 (
	.dataa(!data_out_3),
	.datab(!W_alu_result_3),
	.datac(!W_alu_result_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[3]~3 .extended_lut = "off";
defparam \readdata[3]~3 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \readdata[4]~4 (
	.dataa(!data_out_4),
	.datab(!W_alu_result_3),
	.datac(!W_alu_result_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[4]~4 .extended_lut = "off";
defparam \readdata[4]~4 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \readdata[5]~5 (
	.dataa(!data_out_5),
	.datab(!W_alu_result_3),
	.datac(!W_alu_result_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[5]~5 .extended_lut = "off";
defparam \readdata[5]~5 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!rst1),
	.datab(!wait_latency_counter_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~1 (
	.dataa(!wait_latency_counter_0),
	.datab(!d_write),
	.datac(!write_accepted),
	.datad(!W_alu_result_3),
	.datae(!W_alu_result_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~1 .extended_lut = "off";
defparam \always0~1 .lut_mask = 64'hFFFFFFFBFFFFFFFB;
defparam \always0~1 .shared_arith = "off";

cyclonev_lcell_comb \always0~2 (
	.dataa(!mem_used_1),
	.datab(!W_alu_result_4),
	.datac(!Equal2),
	.datad(!Equal21),
	.datae(!\always0~0_combout ),
	.dataf(!\always0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~2 .extended_lut = "off";
defparam \always0~2 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \always0~2 .shared_arith = "off";

endmodule
