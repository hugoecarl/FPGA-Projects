
module niosLab2 (
	clk_clk,
	leds_export,
	reset_reset_n);	

	input		clk_clk;
	output	[5:0]	leds_export;
	input		reset_reset_n;
endmodule
